magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 3656 4140
<< locali >>
rect 0 0 3656 112
rect 0 0 3656 112
rect 0 0 112 4140
rect 0 4028 3656 4140
rect 3544 0 3656 4140
rect 0 0 3656 112
rect 2746 3390 3070 3610
rect 586 3390 910 3610
<< ptapc >>
rect 28 0 108 80
rect 108 0 188 80
rect 188 0 268 80
rect 268 0 348 80
rect 348 0 428 80
rect 428 0 508 80
rect 508 0 588 80
rect 588 0 668 80
rect 668 0 748 80
rect 748 0 828 80
rect 828 0 908 80
rect 908 0 988 80
rect 988 0 1068 80
rect 1068 0 1148 80
rect 1148 0 1228 80
rect 1228 0 1308 80
rect 1308 0 1388 80
rect 1388 0 1468 80
rect 1468 0 1548 80
rect 1548 0 1628 80
rect 1628 0 1708 80
rect 1708 0 1788 80
rect 1788 0 1868 80
rect 1868 0 1948 80
rect 1948 0 2028 80
rect 2028 0 2108 80
rect 2108 0 2188 80
rect 2188 0 2268 80
rect 2268 0 2348 80
rect 2348 0 2428 80
rect 2428 0 2508 80
rect 2508 0 2588 80
rect 2588 0 2668 80
rect 2668 0 2748 80
rect 2748 0 2828 80
rect 2828 0 2908 80
rect 2908 0 2988 80
rect 2988 0 3068 80
rect 3068 0 3148 80
rect 3148 0 3228 80
rect 3228 0 3308 80
rect 3308 0 3388 80
rect 3388 0 3468 80
rect 3468 0 3548 80
rect 3548 0 3628 80
rect 0 30 80 110
rect 0 110 80 190
rect 0 190 80 270
rect 0 270 80 350
rect 0 350 80 430
rect 0 430 80 510
rect 0 510 80 590
rect 0 590 80 670
rect 0 670 80 750
rect 0 750 80 830
rect 0 830 80 910
rect 0 910 80 990
rect 0 990 80 1070
rect 0 1070 80 1150
rect 0 1150 80 1230
rect 0 1230 80 1310
rect 0 1310 80 1390
rect 0 1390 80 1470
rect 0 1470 80 1550
rect 0 1550 80 1630
rect 0 1630 80 1710
rect 0 1710 80 1790
rect 0 1790 80 1870
rect 0 1870 80 1950
rect 0 1950 80 2030
rect 0 2030 80 2110
rect 0 2110 80 2190
rect 0 2190 80 2270
rect 0 2270 80 2350
rect 0 2350 80 2430
rect 0 2430 80 2510
rect 0 2510 80 2590
rect 0 2590 80 2670
rect 0 2670 80 2750
rect 0 2750 80 2830
rect 0 2830 80 2910
rect 0 2910 80 2990
rect 0 2990 80 3070
rect 0 3070 80 3150
rect 0 3150 80 3230
rect 0 3230 80 3310
rect 0 3310 80 3390
rect 0 3390 80 3470
rect 0 3470 80 3550
rect 0 3550 80 3630
rect 0 3630 80 3710
rect 0 3710 80 3790
rect 0 3790 80 3870
rect 0 3870 80 3950
rect 0 3950 80 4030
rect 0 4030 80 4110
rect 28 4028 108 4108
rect 108 4028 188 4108
rect 188 4028 268 4108
rect 268 4028 348 4108
rect 348 4028 428 4108
rect 428 4028 508 4108
rect 508 4028 588 4108
rect 588 4028 668 4108
rect 668 4028 748 4108
rect 748 4028 828 4108
rect 828 4028 908 4108
rect 908 4028 988 4108
rect 988 4028 1068 4108
rect 1068 4028 1148 4108
rect 1148 4028 1228 4108
rect 1228 4028 1308 4108
rect 1308 4028 1388 4108
rect 1388 4028 1468 4108
rect 1468 4028 1548 4108
rect 1548 4028 1628 4108
rect 1628 4028 1708 4108
rect 1708 4028 1788 4108
rect 1788 4028 1868 4108
rect 1868 4028 1948 4108
rect 1948 4028 2028 4108
rect 2028 4028 2108 4108
rect 2108 4028 2188 4108
rect 2188 4028 2268 4108
rect 2268 4028 2348 4108
rect 2348 4028 2428 4108
rect 2428 4028 2508 4108
rect 2508 4028 2588 4108
rect 2588 4028 2668 4108
rect 2668 4028 2748 4108
rect 2748 4028 2828 4108
rect 2828 4028 2908 4108
rect 2908 4028 2988 4108
rect 2988 4028 3068 4108
rect 3068 4028 3148 4108
rect 3148 4028 3228 4108
rect 3228 4028 3308 4108
rect 3308 4028 3388 4108
rect 3388 4028 3468 4108
rect 3468 4028 3548 4108
rect 3548 4028 3628 4108
rect 3544 30 3624 110
rect 3544 110 3624 190
rect 3544 190 3624 270
rect 3544 270 3624 350
rect 3544 350 3624 430
rect 3544 430 3624 510
rect 3544 510 3624 590
rect 3544 590 3624 670
rect 3544 670 3624 750
rect 3544 750 3624 830
rect 3544 830 3624 910
rect 3544 910 3624 990
rect 3544 990 3624 1070
rect 3544 1070 3624 1150
rect 3544 1150 3624 1230
rect 3544 1230 3624 1310
rect 3544 1310 3624 1390
rect 3544 1390 3624 1470
rect 3544 1470 3624 1550
rect 3544 1550 3624 1630
rect 3544 1630 3624 1710
rect 3544 1710 3624 1790
rect 3544 1790 3624 1870
rect 3544 1870 3624 1950
rect 3544 1950 3624 2030
rect 3544 2030 3624 2110
rect 3544 2110 3624 2190
rect 3544 2190 3624 2270
rect 3544 2270 3624 2350
rect 3544 2350 3624 2430
rect 3544 2430 3624 2510
rect 3544 2510 3624 2590
rect 3544 2590 3624 2670
rect 3544 2670 3624 2750
rect 3544 2750 3624 2830
rect 3544 2830 3624 2910
rect 3544 2910 3624 2990
rect 3544 2990 3624 3070
rect 3544 3070 3624 3150
rect 3544 3150 3624 3230
rect 3544 3230 3624 3310
rect 3544 3310 3624 3390
rect 3544 3390 3624 3470
rect 3544 3470 3624 3550
rect 3544 3550 3624 3630
rect 3544 3630 3624 3710
rect 3544 3710 3624 3790
rect 3544 3790 3624 3870
rect 3544 3870 3624 3950
rect 3544 3950 3624 4030
rect 3544 4030 3624 4110
<< ptap >>
rect 0 0 3656 112
rect 0 0 112 4140
rect 0 4028 3656 4140
rect 3544 0 3656 4140
use SUNTR_RES100 XA1
transform 1 0 640 0 1 640
box 640 640 3016 3500
<< labels >>
flabel locali s 0 0 3656 112 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 2746 3390 3070 3610 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 586 3390 910 3610 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
