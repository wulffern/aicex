magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 11940 4800
<< m1 >>
rect 2490 1810 2850 1870
rect 2580 530 2734 590
rect 2734 770 2940 830
rect 2734 530 2794 838
rect 360 2370 514 2430
rect 514 3090 1920 3150
rect 514 2370 574 3158
rect 1560 2050 1714 2110
rect 1714 2480 2580 2540
rect 1714 2050 1774 2552
rect 720 690 874 750
rect 874 1490 1920 1550
rect 874 690 934 1558
<< locali >>
rect 506 50 720 110
rect 506 370 720 430
rect 506 690 720 750
rect 506 1010 720 1070
rect 506 1330 720 1390
rect 506 1650 720 1710
rect 506 1970 720 2030
rect 506 2290 720 2350
rect 506 50 566 2350
rect 330 130 390 1150
rect 330 1410 390 2430
rect 720 210 874 270
rect 720 530 874 590
rect 720 850 874 910
rect 720 1170 874 1230
rect 874 210 934 1230
rect 720 1490 874 1550
rect 720 1810 874 1870
rect 720 2130 874 2190
rect 720 2450 874 2510
rect 874 1490 934 2510
rect 1470 450 1650 510
rect 2850 770 3030 830
rect 630 1170 810 1230
rect 630 2450 810 2510
<< m2 >>
rect 1560 1730 1714 1798
rect 1714 560 1920 628
rect 1714 560 1782 1798
rect 1154 2130 1920 2198
rect 360 770 1154 838
rect 1154 770 1222 2198
rect 2580 1330 2734 1398
rect 2734 -40 3662 28
rect 2734 -40 2802 1398
<< m3 >>
rect 3438 2680 7740 2748
rect 2942 1810 3438 1878
rect 3438 1810 3506 2748
rect 626 46 810 114
rect 1274 3086 1458 3154
rect 2490 0 2674 4800
rect 1830 0 2014 4800
rect 2490 0 2674 4800
rect 1830 0 2014 4800
use NCHDLR M1
transform 1 0 0 0 1 0
box 0 0 1200 320
use NCHDLR M2
transform 1 0 0 0 1 320
box 0 320 1200 640
use NCHDLR M3
transform 1 0 0 0 1 640
box 0 640 1200 960
use NCHDLR M4
transform 1 0 0 0 1 960
box 0 960 1200 1280
use NCHDLR M5
transform 1 0 0 0 1 1280
box 0 1280 1200 1600
use NCHDLR M6
transform 1 0 0 0 1 1600
box 0 1600 1200 1920
use NCHDLR M7
transform 1 0 0 0 1 1920
box 0 1920 1200 2240
use NCHDLR M8
transform 1 0 0 0 1 2240
box 0 2240 1200 2560
use TAPCELLB_CV XA5b
transform 1 0 1200 0 1 0
box 1200 0 3300 320
use IVX1_CV XA0
transform 1 0 1200 0 1 320
box 1200 320 3300 640
use TGPD_CV XA3
transform 1 0 1200 0 1 640
box 1200 640 3300 1600
use SARBSSWCTRL_CV XA4
transform 1 0 1200 0 1 1600
box 1200 1600 3300 2240
use TIEH_CV XA1
transform 1 0 1200 0 1 2240
box 1200 2240 3300 2560
use TAPCELLB_CV XA7
transform 1 0 1200 0 1 2560
box 1200 2560 3300 2880
use TIEL_CV XA2
transform 1 0 1200 0 1 2880
box 1200 2880 3300 3200
use TAPCELLB_CV XA5
transform 1 0 1200 0 1 3200
box 1200 3200 3300 3520
use CAP_BSSW5_CV XCAPB1
transform 1 0 3480 0 1 0
box 3480 0 11940 4800
use cut_M1M2_2x1 
transform 1 0 2490 0 1 1810
box 2490 1810 2674 1878
use cut_M2M4_2x1 
transform 1 0 2850 0 1 1810
box 2850 1810 3034 1878
use cut_M1M2_2x1 
transform 1 0 2490 0 1 530
box 2490 530 2674 598
use cut_M1M2_2x1 
transform 1 0 2850 0 1 770
box 2850 770 3034 838
use cut_M1M3_2x1 
transform 1 0 1470 0 1 1730
box 1470 1730 1654 1798
use cut_M1M3_2x1 
transform 1 0 1830 0 1 564
box 1830 564 2014 632
use cut_M1M2_2x1 
transform 1 0 270 0 1 2370
box 270 2370 454 2438
use cut_M1M2_2x1 
transform 1 0 1830 0 1 3090
box 1830 3090 2014 3158
use cut_M1M2_2x1 
transform 1 0 1470 0 1 2050
box 1470 2050 1654 2118
use cut_M1M2_2x1 
transform 1 0 2490 0 1 2484
box 2490 2484 2674 2552
use cut_M1M2_2x1 
transform 1 0 630 0 1 690
box 630 690 814 758
use cut_M1M2_2x1 
transform 1 0 1830 0 1 1490
box 1830 1490 2014 1558
use cut_M1M3_2x1 
transform 1 0 1826 0 1 2130
box 1826 2130 2010 2198
use cut_M1M3_2x1 
transform 1 0 266 0 1 770
box 266 770 450 838
use cut_M1M3_2x1 
transform 1 0 2490 0 1 1330
box 2490 1330 2674 1398
use cut_M3M4_2x1 
transform 1 0 3570 0 1 -40
box 3570 -40 3754 28
use cut_M1M4_2x1 
transform 1 0 626 0 1 46
box 626 46 810 114
use cut_M2M4_2x1 
transform 1 0 1274 0 1 3086
box 1274 3086 1458 3154
<< labels >>
flabel m3 s 626 46 810 114 0 FreeSans 400 0 0 0 VI
port 1 nsew
flabel m3 s 1274 3086 1458 3154 0 FreeSans 400 0 0 0 TIE_L
port 2 nsew
flabel locali s 1470 450 1650 510 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel locali s 2850 770 3030 830 0 FreeSans 400 0 0 0 CKN
port 4 nsew
flabel locali s 630 1170 810 1230 0 FreeSans 400 0 0 0 VO1
port 5 nsew
flabel locali s 630 2450 810 2510 0 FreeSans 400 0 0 0 VO2
port 6 nsew
flabel m3 s 2490 0 2674 4800 0 FreeSans 400 0 0 0 AVDD
port 7 nsew
flabel m3 s 1830 0 2014 4800 0 FreeSans 400 0 0 0 AVSS
port 8 nsew
<< end >>
