magic
tech sky130A
magscale 1 2
timestamp 1660740729
<< checkpaint >>
rect 0 0 1440 352
<< ndiff >>
rect 756 220 972 308
rect 756 132 972 220
rect 756 44 972 132
<< ptap >>
rect -108 308 108 396
rect -108 220 108 308
rect -108 132 108 220
rect -108 44 108 132
rect -108 -44 108 44
<< poly >>
rect 324 334 1044 370
rect 324 158 1044 194
rect 324 -18 1044 18
rect 324 132 540 220
<< locali >>
rect 324 146 540 206
rect -108 308 108 396
rect -108 220 108 308
rect 756 234 972 294
rect 756 234 972 294
rect -108 132 108 220
rect -108 132 108 220
rect 324 146 540 206
rect -108 44 108 132
rect 756 58 972 118
rect 756 58 972 118
rect -108 -44 108 44
<< pcontact >>
rect 348 176 396 198
rect 348 154 396 176
rect 396 176 468 198
rect 396 154 468 176
rect 468 176 516 198
rect 468 154 516 176
<< ptapc >>
rect -36 220 36 308
rect -36 44 36 132
<< ndcontact >>
rect 780 264 828 286
rect 780 242 828 264
rect 828 264 900 286
rect 828 242 900 264
rect 900 264 948 286
rect 900 242 948 264
rect 780 88 828 110
rect 780 66 828 88
rect 828 88 900 110
rect 828 66 900 88
rect 900 88 948 110
rect 900 66 948 88
<< pwell >>
rect -180 -132 1260 484
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 756 234 972 294 0 FreeSans 400 0 0 0 S
port 3 nsew
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 756 58 972 118 0 FreeSans 400 0 0 0 D
port 1 nsew
<< end >>
