magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 960
<< locali >>
rect 720 850 874 910
rect 874 850 1380 910
rect 874 850 934 910
rect 1710 130 1770 830
rect 690 210 750 430
rect 690 530 750 750
rect 1350 210 1410 430
rect 1350 530 1410 750
rect 2010 120 2190 200
rect -90 120 90 200
rect 270 130 450 190
rect 1650 770 1830 830
rect 270 770 450 830
rect 270 450 450 510
rect 630 850 810 910
<< m3 >>
rect 1290 0 1474 960
rect 630 0 814 960
rect 1290 0 1474 960
rect 630 0 814 960
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1050 960
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL MP2
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use cut_M1M4_2x1 
transform 1 0 1290 0 1 50
box 1290 50 1474 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
<< labels >>
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel locali s 1650 770 1830 830 0 FreeSans 400 0 0 0 RST_N
port 4 nsew
flabel locali s 270 770 450 830 0 FreeSans 400 0 0 0 EN
port 5 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 LCK_N
port 6 nsew
flabel locali s 630 850 810 910 0 FreeSans 400 0 0 0 CHL
port 7 nsew
flabel m3 s 1290 0 1474 960 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 960 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
