magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 116 0 11404 11964
<< m1 >>
rect 2188 4596 2248 11904
rect 2188 4596 2248 11904
rect 2000 132 2060 11904
rect 2000 132 2060 11904
rect 1812 9060 1872 11904
rect 1812 9060 1872 11904
rect 1624 1620 1684 11904
rect 1624 1620 1684 11904
rect 1436 3328 1496 11904
rect 1436 3328 1496 11904
rect 1248 7792 1308 11904
rect 1248 7792 1308 11904
rect 1060 7572 1120 11904
rect 1060 7572 1120 11904
rect 872 8232 932 11904
rect 872 8232 932 11904
rect 684 3768 744 11904
rect 684 3768 744 11904
rect 496 3988 556 11904
rect 496 3988 556 11904
rect 308 3548 368 11904
rect 308 3548 368 11904
rect 120 4208 180 11904
rect 120 4208 180 11904
rect 2756 0 11336 68
<< m2 >>
rect 2444 4654 2248 4722
rect 2444 5754 2248 5822
rect 2444 5094 2248 5162
rect 2444 5534 2248 5602
rect 2444 5314 2248 5382
rect 2444 4874 2248 4942
rect 2444 4654 2248 4722
rect 2444 5754 2248 5822
rect 2444 5094 2248 5162
rect 2444 5534 2248 5602
rect 2444 5314 2248 5382
rect 2444 4874 2248 4942
rect 2444 4654 2248 4722
rect 2444 5754 2248 5822
rect 2444 5094 2248 5162
rect 2444 5534 2248 5602
rect 2444 5314 2248 5382
rect 2444 4874 2248 4942
rect 2444 4654 2248 4722
rect 2444 5754 2248 5822
rect 2444 5094 2248 5162
rect 2444 5534 2248 5602
rect 2444 5314 2248 5382
rect 2444 4874 2248 4942
rect 2444 4654 2248 4722
rect 2444 5754 2248 5822
rect 2444 5094 2248 5162
rect 2444 5534 2248 5602
rect 2444 5314 2248 5382
rect 2444 4874 2248 4942
rect 2444 4654 2248 4722
rect 2444 5754 2248 5822
rect 2444 5094 2248 5162
rect 2444 5534 2248 5602
rect 2444 5314 2248 5382
rect 2444 4874 2248 4942
rect 2444 10606 2248 10674
rect 2444 11706 2248 11774
rect 2444 11046 2248 11114
rect 2444 11486 2248 11554
rect 2444 11266 2248 11334
rect 2444 10826 2248 10894
rect 2444 10606 2248 10674
rect 2444 11706 2248 11774
rect 2444 11046 2248 11114
rect 2444 11486 2248 11554
rect 2444 11266 2248 11334
rect 2444 10826 2248 10894
rect 2444 10606 2248 10674
rect 2444 11706 2248 11774
rect 2444 11046 2248 11114
rect 2444 11486 2248 11554
rect 2444 11266 2248 11334
rect 2444 10826 2248 10894
rect 2444 10606 2248 10674
rect 2444 11706 2248 11774
rect 2444 11046 2248 11114
rect 2444 11486 2248 11554
rect 2444 11266 2248 11334
rect 2444 10826 2248 10894
rect 2444 10606 2248 10674
rect 2444 11706 2248 11774
rect 2444 11046 2248 11114
rect 2444 11486 2248 11554
rect 2444 11266 2248 11334
rect 2444 10826 2248 10894
rect 2444 10606 2248 10674
rect 2444 11706 2248 11774
rect 2444 11046 2248 11114
rect 2444 11486 2248 11554
rect 2444 11266 2248 11334
rect 2444 10826 2248 10894
rect 2444 190 2060 258
rect 2444 1290 2060 1358
rect 2444 630 2060 698
rect 2444 1070 2060 1138
rect 2444 850 2060 918
rect 2444 410 2060 478
rect 2444 190 2060 258
rect 2444 1290 2060 1358
rect 2444 630 2060 698
rect 2444 1070 2060 1138
rect 2444 850 2060 918
rect 2444 410 2060 478
rect 2444 190 2060 258
rect 2444 1290 2060 1358
rect 2444 630 2060 698
rect 2444 1070 2060 1138
rect 2444 850 2060 918
rect 2444 410 2060 478
rect 2444 190 2060 258
rect 2444 1290 2060 1358
rect 2444 630 2060 698
rect 2444 1070 2060 1138
rect 2444 850 2060 918
rect 2444 410 2060 478
rect 2444 190 2060 258
rect 2444 1290 2060 1358
rect 2444 630 2060 698
rect 2444 1070 2060 1138
rect 2444 850 2060 918
rect 2444 410 2060 478
rect 2444 190 2060 258
rect 2444 1290 2060 1358
rect 2444 630 2060 698
rect 2444 1070 2060 1138
rect 2444 850 2060 918
rect 2444 410 2060 478
rect 2444 6142 2060 6210
rect 2444 7242 2060 7310
rect 2444 6582 2060 6650
rect 2444 7022 2060 7090
rect 2444 6802 2060 6870
rect 2444 6362 2060 6430
rect 2444 6142 2060 6210
rect 2444 7242 2060 7310
rect 2444 6582 2060 6650
rect 2444 7022 2060 7090
rect 2444 6802 2060 6870
rect 2444 6362 2060 6430
rect 2444 6142 2060 6210
rect 2444 7242 2060 7310
rect 2444 6582 2060 6650
rect 2444 7022 2060 7090
rect 2444 6802 2060 6870
rect 2444 6362 2060 6430
rect 2444 6142 2060 6210
rect 2444 7242 2060 7310
rect 2444 6582 2060 6650
rect 2444 7022 2060 7090
rect 2444 6802 2060 6870
rect 2444 6362 2060 6430
rect 2444 6142 2060 6210
rect 2444 7242 2060 7310
rect 2444 6582 2060 6650
rect 2444 7022 2060 7090
rect 2444 6802 2060 6870
rect 2444 6362 2060 6430
rect 2444 6142 2060 6210
rect 2444 7242 2060 7310
rect 2444 6582 2060 6650
rect 2444 7022 2060 7090
rect 2444 6802 2060 6870
rect 2444 6362 2060 6430
rect 2444 9118 1872 9186
rect 2444 10218 1872 10286
rect 2444 9558 1872 9626
rect 2444 9998 1872 10066
rect 2444 9778 1872 9846
rect 2444 9338 1872 9406
rect 2444 9118 1872 9186
rect 2444 10218 1872 10286
rect 2444 9558 1872 9626
rect 2444 9998 1872 10066
rect 2444 9778 1872 9846
rect 2444 9338 1872 9406
rect 2444 9118 1872 9186
rect 2444 10218 1872 10286
rect 2444 9558 1872 9626
rect 2444 9998 1872 10066
rect 2444 9778 1872 9846
rect 2444 9338 1872 9406
rect 2444 9118 1872 9186
rect 2444 10218 1872 10286
rect 2444 9558 1872 9626
rect 2444 9998 1872 10066
rect 2444 9778 1872 9846
rect 2444 9338 1872 9406
rect 2444 9118 1872 9186
rect 2444 10218 1872 10286
rect 2444 9558 1872 9626
rect 2444 9998 1872 10066
rect 2444 9778 1872 9846
rect 2444 9338 1872 9406
rect 2444 9118 1872 9186
rect 2444 10218 1872 10286
rect 2444 9558 1872 9626
rect 2444 9998 1872 10066
rect 2444 9778 1872 9846
rect 2444 9338 1872 9406
rect 2444 1678 1684 1746
rect 2444 2778 1684 2846
rect 2444 2118 1684 2186
rect 2444 2558 1684 2626
rect 2444 2338 1684 2406
rect 2444 1898 1684 1966
rect 2444 1678 1684 1746
rect 2444 2778 1684 2846
rect 2444 2118 1684 2186
rect 2444 2558 1684 2626
rect 2444 2338 1684 2406
rect 2444 1898 1684 1966
rect 2444 1678 1684 1746
rect 2444 2778 1684 2846
rect 2444 2118 1684 2186
rect 2444 2558 1684 2626
rect 2444 2338 1684 2406
rect 2444 1898 1684 1966
rect 2444 1678 1684 1746
rect 2444 2778 1684 2846
rect 2444 2118 1684 2186
rect 2444 2558 1684 2626
rect 2444 2338 1684 2406
rect 2444 1898 1684 1966
rect 2444 1678 1684 1746
rect 2444 2778 1684 2846
rect 2444 2118 1684 2186
rect 2444 2558 1684 2626
rect 2444 2338 1684 2406
rect 2444 1898 1684 1966
rect 2444 1678 1684 1746
rect 2444 2778 1684 2846
rect 2444 2118 1684 2186
rect 2444 2558 1684 2626
rect 2444 2338 1684 2406
rect 2444 1898 1684 1966
rect 2444 3386 1496 3454
rect 2444 7850 1308 7918
rect 2444 7630 1120 7698
rect 2444 8730 1120 8798
rect 2444 8070 1120 8138
rect 2444 8510 1120 8578
rect 2444 7630 1120 7698
rect 2444 8730 1120 8798
rect 2444 8070 1120 8138
rect 2444 8510 1120 8578
rect 2444 7630 1120 7698
rect 2444 8730 1120 8798
rect 2444 8070 1120 8138
rect 2444 8510 1120 8578
rect 2444 7630 1120 7698
rect 2444 8730 1120 8798
rect 2444 8070 1120 8138
rect 2444 8510 1120 8578
rect 2444 8290 932 8358
rect 2444 3826 744 3894
rect 2444 4046 556 4114
rect 2444 3606 368 3674
rect 2444 4266 180 4334
<< m3 >>
rect 2756 10416 2824 11964
use CAP32C_CV XC1
transform 1 0 2444 0 1 0
box 2444 0 11404 1488
use CAP32C_CV XC64a<0>
transform 1 0 2444 0 1 1488
box 2444 1488 11404 2976
use CAP32C_CV XC32a<0>
transform 1 0 2444 0 1 2976
box 2444 2976 11404 4464
use CAP32C_CV XC128a<1>
transform 1 0 2444 0 1 4464
box 2444 4464 11404 5952
use CAP32C_CV XC128b<2>
transform 1 0 2444 0 1 5952
box 2444 5952 11404 7440
use CAP32C_CV X16ab
transform 1 0 2444 0 1 7440
box 2444 7440 11404 8928
use CAP32C_CV XC64b<1>
transform 1 0 2444 0 1 8928
box 2444 8928 11404 10416
use CAP32C_CV XC0
transform 1 0 2444 0 1 10416
box 2444 10416 11404 11904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4654
box 2444 4654 2628 4722
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4596
box 2184 4596 2252 4780
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5754
box 2444 5754 2628 5822
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5696
box 2184 5696 2252 5880
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5094
box 2444 5094 2628 5162
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5036
box 2184 5036 2252 5220
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5534
box 2444 5534 2628 5602
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5476
box 2184 5476 2252 5660
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5314
box 2444 5314 2628 5382
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5256
box 2184 5256 2252 5440
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4874
box 2444 4874 2628 4942
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4816
box 2184 4816 2252 5000
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4654
box 2444 4654 2628 4722
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4596
box 2184 4596 2252 4780
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5754
box 2444 5754 2628 5822
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5696
box 2184 5696 2252 5880
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5094
box 2444 5094 2628 5162
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5036
box 2184 5036 2252 5220
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5534
box 2444 5534 2628 5602
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5476
box 2184 5476 2252 5660
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5314
box 2444 5314 2628 5382
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5256
box 2184 5256 2252 5440
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4874
box 2444 4874 2628 4942
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4816
box 2184 4816 2252 5000
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4654
box 2444 4654 2628 4722
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4596
box 2184 4596 2252 4780
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5754
box 2444 5754 2628 5822
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5696
box 2184 5696 2252 5880
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5094
box 2444 5094 2628 5162
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5036
box 2184 5036 2252 5220
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5534
box 2444 5534 2628 5602
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5476
box 2184 5476 2252 5660
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5314
box 2444 5314 2628 5382
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5256
box 2184 5256 2252 5440
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4874
box 2444 4874 2628 4942
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4816
box 2184 4816 2252 5000
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4654
box 2444 4654 2628 4722
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4596
box 2184 4596 2252 4780
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5754
box 2444 5754 2628 5822
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5696
box 2184 5696 2252 5880
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5094
box 2444 5094 2628 5162
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5036
box 2184 5036 2252 5220
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5534
box 2444 5534 2628 5602
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5476
box 2184 5476 2252 5660
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5314
box 2444 5314 2628 5382
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5256
box 2184 5256 2252 5440
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4874
box 2444 4874 2628 4942
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4816
box 2184 4816 2252 5000
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4654
box 2444 4654 2628 4722
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4596
box 2184 4596 2252 4780
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5754
box 2444 5754 2628 5822
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5696
box 2184 5696 2252 5880
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5094
box 2444 5094 2628 5162
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5036
box 2184 5036 2252 5220
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5534
box 2444 5534 2628 5602
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5476
box 2184 5476 2252 5660
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5314
box 2444 5314 2628 5382
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5256
box 2184 5256 2252 5440
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4874
box 2444 4874 2628 4942
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4816
box 2184 4816 2252 5000
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4654
box 2444 4654 2628 4722
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4596
box 2184 4596 2252 4780
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5754
box 2444 5754 2628 5822
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5696
box 2184 5696 2252 5880
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5094
box 2444 5094 2628 5162
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5036
box 2184 5036 2252 5220
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5534
box 2444 5534 2628 5602
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5476
box 2184 5476 2252 5660
use cut_M1M3_2x1 
transform 1 0 2444 0 1 5314
box 2444 5314 2628 5382
use cut_M2M3_1x2 
transform 1 0 2184 0 1 5256
box 2184 5256 2252 5440
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4874
box 2444 4874 2628 4942
use cut_M2M3_1x2 
transform 1 0 2184 0 1 4816
box 2184 4816 2252 5000
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10606
box 2444 10606 2628 10674
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10548
box 2184 10548 2252 10732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11706
box 2444 11706 2628 11774
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11648
box 2184 11648 2252 11832
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11046
box 2444 11046 2628 11114
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10988
box 2184 10988 2252 11172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11486
box 2444 11486 2628 11554
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11428
box 2184 11428 2252 11612
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11266
box 2444 11266 2628 11334
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11208
box 2184 11208 2252 11392
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10826
box 2444 10826 2628 10894
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10768
box 2184 10768 2252 10952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10606
box 2444 10606 2628 10674
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10548
box 2184 10548 2252 10732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11706
box 2444 11706 2628 11774
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11648
box 2184 11648 2252 11832
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11046
box 2444 11046 2628 11114
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10988
box 2184 10988 2252 11172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11486
box 2444 11486 2628 11554
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11428
box 2184 11428 2252 11612
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11266
box 2444 11266 2628 11334
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11208
box 2184 11208 2252 11392
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10826
box 2444 10826 2628 10894
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10768
box 2184 10768 2252 10952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10606
box 2444 10606 2628 10674
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10548
box 2184 10548 2252 10732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11706
box 2444 11706 2628 11774
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11648
box 2184 11648 2252 11832
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11046
box 2444 11046 2628 11114
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10988
box 2184 10988 2252 11172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11486
box 2444 11486 2628 11554
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11428
box 2184 11428 2252 11612
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11266
box 2444 11266 2628 11334
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11208
box 2184 11208 2252 11392
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10826
box 2444 10826 2628 10894
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10768
box 2184 10768 2252 10952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10606
box 2444 10606 2628 10674
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10548
box 2184 10548 2252 10732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11706
box 2444 11706 2628 11774
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11648
box 2184 11648 2252 11832
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11046
box 2444 11046 2628 11114
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10988
box 2184 10988 2252 11172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11486
box 2444 11486 2628 11554
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11428
box 2184 11428 2252 11612
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11266
box 2444 11266 2628 11334
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11208
box 2184 11208 2252 11392
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10826
box 2444 10826 2628 10894
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10768
box 2184 10768 2252 10952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10606
box 2444 10606 2628 10674
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10548
box 2184 10548 2252 10732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11706
box 2444 11706 2628 11774
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11648
box 2184 11648 2252 11832
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11046
box 2444 11046 2628 11114
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10988
box 2184 10988 2252 11172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11486
box 2444 11486 2628 11554
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11428
box 2184 11428 2252 11612
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11266
box 2444 11266 2628 11334
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11208
box 2184 11208 2252 11392
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10826
box 2444 10826 2628 10894
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10768
box 2184 10768 2252 10952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10606
box 2444 10606 2628 10674
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10548
box 2184 10548 2252 10732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11706
box 2444 11706 2628 11774
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11648
box 2184 11648 2252 11832
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11046
box 2444 11046 2628 11114
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10988
box 2184 10988 2252 11172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11486
box 2444 11486 2628 11554
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11428
box 2184 11428 2252 11612
use cut_M1M3_2x1 
transform 1 0 2444 0 1 11266
box 2444 11266 2628 11334
use cut_M2M3_1x2 
transform 1 0 2184 0 1 11208
box 2184 11208 2252 11392
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10826
box 2444 10826 2628 10894
use cut_M2M3_1x2 
transform 1 0 2184 0 1 10768
box 2184 10768 2252 10952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use cut_M2M3_1x2 
transform 1 0 1996 0 1 132
box 1996 132 2064 316
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1290
box 2444 1290 2628 1358
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1232
box 1996 1232 2064 1416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 630
box 2444 630 2628 698
use cut_M2M3_1x2 
transform 1 0 1996 0 1 572
box 1996 572 2064 756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1070
box 2444 1070 2628 1138
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1012
box 1996 1012 2064 1196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 850
box 2444 850 2628 918
use cut_M2M3_1x2 
transform 1 0 1996 0 1 792
box 1996 792 2064 976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 410
box 2444 410 2628 478
use cut_M2M3_1x2 
transform 1 0 1996 0 1 352
box 1996 352 2064 536
use cut_M1M3_2x1 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use cut_M2M3_1x2 
transform 1 0 1996 0 1 132
box 1996 132 2064 316
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1290
box 2444 1290 2628 1358
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1232
box 1996 1232 2064 1416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 630
box 2444 630 2628 698
use cut_M2M3_1x2 
transform 1 0 1996 0 1 572
box 1996 572 2064 756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1070
box 2444 1070 2628 1138
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1012
box 1996 1012 2064 1196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 850
box 2444 850 2628 918
use cut_M2M3_1x2 
transform 1 0 1996 0 1 792
box 1996 792 2064 976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 410
box 2444 410 2628 478
use cut_M2M3_1x2 
transform 1 0 1996 0 1 352
box 1996 352 2064 536
use cut_M1M3_2x1 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use cut_M2M3_1x2 
transform 1 0 1996 0 1 132
box 1996 132 2064 316
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1290
box 2444 1290 2628 1358
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1232
box 1996 1232 2064 1416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 630
box 2444 630 2628 698
use cut_M2M3_1x2 
transform 1 0 1996 0 1 572
box 1996 572 2064 756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1070
box 2444 1070 2628 1138
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1012
box 1996 1012 2064 1196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 850
box 2444 850 2628 918
use cut_M2M3_1x2 
transform 1 0 1996 0 1 792
box 1996 792 2064 976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 410
box 2444 410 2628 478
use cut_M2M3_1x2 
transform 1 0 1996 0 1 352
box 1996 352 2064 536
use cut_M1M3_2x1 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use cut_M2M3_1x2 
transform 1 0 1996 0 1 132
box 1996 132 2064 316
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1290
box 2444 1290 2628 1358
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1232
box 1996 1232 2064 1416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 630
box 2444 630 2628 698
use cut_M2M3_1x2 
transform 1 0 1996 0 1 572
box 1996 572 2064 756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1070
box 2444 1070 2628 1138
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1012
box 1996 1012 2064 1196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 850
box 2444 850 2628 918
use cut_M2M3_1x2 
transform 1 0 1996 0 1 792
box 1996 792 2064 976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 410
box 2444 410 2628 478
use cut_M2M3_1x2 
transform 1 0 1996 0 1 352
box 1996 352 2064 536
use cut_M1M3_2x1 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use cut_M2M3_1x2 
transform 1 0 1996 0 1 132
box 1996 132 2064 316
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1290
box 2444 1290 2628 1358
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1232
box 1996 1232 2064 1416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 630
box 2444 630 2628 698
use cut_M2M3_1x2 
transform 1 0 1996 0 1 572
box 1996 572 2064 756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1070
box 2444 1070 2628 1138
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1012
box 1996 1012 2064 1196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 850
box 2444 850 2628 918
use cut_M2M3_1x2 
transform 1 0 1996 0 1 792
box 1996 792 2064 976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 410
box 2444 410 2628 478
use cut_M2M3_1x2 
transform 1 0 1996 0 1 352
box 1996 352 2064 536
use cut_M1M3_2x1 
transform 1 0 2444 0 1 190
box 2444 190 2628 258
use cut_M2M3_1x2 
transform 1 0 1996 0 1 132
box 1996 132 2064 316
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1290
box 2444 1290 2628 1358
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1232
box 1996 1232 2064 1416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 630
box 2444 630 2628 698
use cut_M2M3_1x2 
transform 1 0 1996 0 1 572
box 1996 572 2064 756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1070
box 2444 1070 2628 1138
use cut_M2M3_1x2 
transform 1 0 1996 0 1 1012
box 1996 1012 2064 1196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 850
box 2444 850 2628 918
use cut_M2M3_1x2 
transform 1 0 1996 0 1 792
box 1996 792 2064 976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 410
box 2444 410 2628 478
use cut_M2M3_1x2 
transform 1 0 1996 0 1 352
box 1996 352 2064 536
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6142
box 2444 6142 2628 6210
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6084
box 1996 6084 2064 6268
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7242
box 2444 7242 2628 7310
use cut_M2M3_1x2 
transform 1 0 1996 0 1 7184
box 1996 7184 2064 7368
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6582
box 2444 6582 2628 6650
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6524
box 1996 6524 2064 6708
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7022
box 2444 7022 2628 7090
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6964
box 1996 6964 2064 7148
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6802
box 2444 6802 2628 6870
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6744
box 1996 6744 2064 6928
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6362
box 2444 6362 2628 6430
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6304
box 1996 6304 2064 6488
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6142
box 2444 6142 2628 6210
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6084
box 1996 6084 2064 6268
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7242
box 2444 7242 2628 7310
use cut_M2M3_1x2 
transform 1 0 1996 0 1 7184
box 1996 7184 2064 7368
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6582
box 2444 6582 2628 6650
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6524
box 1996 6524 2064 6708
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7022
box 2444 7022 2628 7090
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6964
box 1996 6964 2064 7148
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6802
box 2444 6802 2628 6870
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6744
box 1996 6744 2064 6928
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6362
box 2444 6362 2628 6430
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6304
box 1996 6304 2064 6488
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6142
box 2444 6142 2628 6210
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6084
box 1996 6084 2064 6268
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7242
box 2444 7242 2628 7310
use cut_M2M3_1x2 
transform 1 0 1996 0 1 7184
box 1996 7184 2064 7368
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6582
box 2444 6582 2628 6650
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6524
box 1996 6524 2064 6708
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7022
box 2444 7022 2628 7090
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6964
box 1996 6964 2064 7148
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6802
box 2444 6802 2628 6870
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6744
box 1996 6744 2064 6928
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6362
box 2444 6362 2628 6430
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6304
box 1996 6304 2064 6488
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6142
box 2444 6142 2628 6210
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6084
box 1996 6084 2064 6268
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7242
box 2444 7242 2628 7310
use cut_M2M3_1x2 
transform 1 0 1996 0 1 7184
box 1996 7184 2064 7368
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6582
box 2444 6582 2628 6650
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6524
box 1996 6524 2064 6708
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7022
box 2444 7022 2628 7090
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6964
box 1996 6964 2064 7148
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6802
box 2444 6802 2628 6870
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6744
box 1996 6744 2064 6928
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6362
box 2444 6362 2628 6430
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6304
box 1996 6304 2064 6488
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6142
box 2444 6142 2628 6210
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6084
box 1996 6084 2064 6268
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7242
box 2444 7242 2628 7310
use cut_M2M3_1x2 
transform 1 0 1996 0 1 7184
box 1996 7184 2064 7368
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6582
box 2444 6582 2628 6650
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6524
box 1996 6524 2064 6708
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7022
box 2444 7022 2628 7090
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6964
box 1996 6964 2064 7148
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6802
box 2444 6802 2628 6870
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6744
box 1996 6744 2064 6928
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6362
box 2444 6362 2628 6430
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6304
box 1996 6304 2064 6488
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6142
box 2444 6142 2628 6210
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6084
box 1996 6084 2064 6268
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7242
box 2444 7242 2628 7310
use cut_M2M3_1x2 
transform 1 0 1996 0 1 7184
box 1996 7184 2064 7368
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6582
box 2444 6582 2628 6650
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6524
box 1996 6524 2064 6708
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7022
box 2444 7022 2628 7090
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6964
box 1996 6964 2064 7148
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6802
box 2444 6802 2628 6870
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6744
box 1996 6744 2064 6928
use cut_M1M3_2x1 
transform 1 0 2444 0 1 6362
box 2444 6362 2628 6430
use cut_M2M3_1x2 
transform 1 0 1996 0 1 6304
box 1996 6304 2064 6488
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9118
box 2444 9118 2628 9186
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9060
box 1808 9060 1876 9244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10218
box 2444 10218 2628 10286
use cut_M2M3_1x2 
transform 1 0 1808 0 1 10160
box 1808 10160 1876 10344
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9558
box 2444 9558 2628 9626
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9500
box 1808 9500 1876 9684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9998
box 2444 9998 2628 10066
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9940
box 1808 9940 1876 10124
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9778
box 2444 9778 2628 9846
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9720
box 1808 9720 1876 9904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9338
box 2444 9338 2628 9406
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9280
box 1808 9280 1876 9464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9118
box 2444 9118 2628 9186
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9060
box 1808 9060 1876 9244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10218
box 2444 10218 2628 10286
use cut_M2M3_1x2 
transform 1 0 1808 0 1 10160
box 1808 10160 1876 10344
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9558
box 2444 9558 2628 9626
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9500
box 1808 9500 1876 9684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9998
box 2444 9998 2628 10066
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9940
box 1808 9940 1876 10124
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9778
box 2444 9778 2628 9846
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9720
box 1808 9720 1876 9904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9338
box 2444 9338 2628 9406
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9280
box 1808 9280 1876 9464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9118
box 2444 9118 2628 9186
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9060
box 1808 9060 1876 9244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10218
box 2444 10218 2628 10286
use cut_M2M3_1x2 
transform 1 0 1808 0 1 10160
box 1808 10160 1876 10344
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9558
box 2444 9558 2628 9626
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9500
box 1808 9500 1876 9684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9998
box 2444 9998 2628 10066
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9940
box 1808 9940 1876 10124
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9778
box 2444 9778 2628 9846
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9720
box 1808 9720 1876 9904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9338
box 2444 9338 2628 9406
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9280
box 1808 9280 1876 9464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9118
box 2444 9118 2628 9186
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9060
box 1808 9060 1876 9244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10218
box 2444 10218 2628 10286
use cut_M2M3_1x2 
transform 1 0 1808 0 1 10160
box 1808 10160 1876 10344
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9558
box 2444 9558 2628 9626
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9500
box 1808 9500 1876 9684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9998
box 2444 9998 2628 10066
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9940
box 1808 9940 1876 10124
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9778
box 2444 9778 2628 9846
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9720
box 1808 9720 1876 9904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9338
box 2444 9338 2628 9406
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9280
box 1808 9280 1876 9464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9118
box 2444 9118 2628 9186
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9060
box 1808 9060 1876 9244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10218
box 2444 10218 2628 10286
use cut_M2M3_1x2 
transform 1 0 1808 0 1 10160
box 1808 10160 1876 10344
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9558
box 2444 9558 2628 9626
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9500
box 1808 9500 1876 9684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9998
box 2444 9998 2628 10066
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9940
box 1808 9940 1876 10124
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9778
box 2444 9778 2628 9846
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9720
box 1808 9720 1876 9904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9338
box 2444 9338 2628 9406
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9280
box 1808 9280 1876 9464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9118
box 2444 9118 2628 9186
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9060
box 1808 9060 1876 9244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 10218
box 2444 10218 2628 10286
use cut_M2M3_1x2 
transform 1 0 1808 0 1 10160
box 1808 10160 1876 10344
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9558
box 2444 9558 2628 9626
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9500
box 1808 9500 1876 9684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9998
box 2444 9998 2628 10066
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9940
box 1808 9940 1876 10124
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9778
box 2444 9778 2628 9846
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9720
box 1808 9720 1876 9904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 9338
box 2444 9338 2628 9406
use cut_M2M3_1x2 
transform 1 0 1808 0 1 9280
box 1808 9280 1876 9464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1678
box 2444 1678 2628 1746
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1620
box 1620 1620 1688 1804
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2778
box 2444 2778 2628 2846
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2720
box 1620 2720 1688 2904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2118
box 2444 2118 2628 2186
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2060
box 1620 2060 1688 2244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2558
box 2444 2558 2628 2626
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2500
box 1620 2500 1688 2684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2338
box 2444 2338 2628 2406
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2280
box 1620 2280 1688 2464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1898
box 2444 1898 2628 1966
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1840
box 1620 1840 1688 2024
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1678
box 2444 1678 2628 1746
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1620
box 1620 1620 1688 1804
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2778
box 2444 2778 2628 2846
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2720
box 1620 2720 1688 2904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2118
box 2444 2118 2628 2186
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2060
box 1620 2060 1688 2244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2558
box 2444 2558 2628 2626
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2500
box 1620 2500 1688 2684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2338
box 2444 2338 2628 2406
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2280
box 1620 2280 1688 2464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1898
box 2444 1898 2628 1966
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1840
box 1620 1840 1688 2024
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1678
box 2444 1678 2628 1746
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1620
box 1620 1620 1688 1804
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2778
box 2444 2778 2628 2846
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2720
box 1620 2720 1688 2904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2118
box 2444 2118 2628 2186
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2060
box 1620 2060 1688 2244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2558
box 2444 2558 2628 2626
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2500
box 1620 2500 1688 2684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2338
box 2444 2338 2628 2406
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2280
box 1620 2280 1688 2464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1898
box 2444 1898 2628 1966
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1840
box 1620 1840 1688 2024
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1678
box 2444 1678 2628 1746
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1620
box 1620 1620 1688 1804
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2778
box 2444 2778 2628 2846
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2720
box 1620 2720 1688 2904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2118
box 2444 2118 2628 2186
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2060
box 1620 2060 1688 2244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2558
box 2444 2558 2628 2626
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2500
box 1620 2500 1688 2684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2338
box 2444 2338 2628 2406
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2280
box 1620 2280 1688 2464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1898
box 2444 1898 2628 1966
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1840
box 1620 1840 1688 2024
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1678
box 2444 1678 2628 1746
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1620
box 1620 1620 1688 1804
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2778
box 2444 2778 2628 2846
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2720
box 1620 2720 1688 2904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2118
box 2444 2118 2628 2186
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2060
box 1620 2060 1688 2244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2558
box 2444 2558 2628 2626
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2500
box 1620 2500 1688 2684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2338
box 2444 2338 2628 2406
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2280
box 1620 2280 1688 2464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1898
box 2444 1898 2628 1966
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1840
box 1620 1840 1688 2024
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1678
box 2444 1678 2628 1746
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1620
box 1620 1620 1688 1804
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2778
box 2444 2778 2628 2846
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2720
box 1620 2720 1688 2904
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2118
box 2444 2118 2628 2186
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2060
box 1620 2060 1688 2244
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2558
box 2444 2558 2628 2626
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2500
box 1620 2500 1688 2684
use cut_M1M3_2x1 
transform 1 0 2444 0 1 2338
box 2444 2338 2628 2406
use cut_M2M3_1x2 
transform 1 0 1620 0 1 2280
box 1620 2280 1688 2464
use cut_M1M3_2x1 
transform 1 0 2444 0 1 1898
box 2444 1898 2628 1966
use cut_M2M3_1x2 
transform 1 0 1620 0 1 1840
box 1620 1840 1688 2024
use cut_M1M3_2x1 
transform 1 0 2444 0 1 3386
box 2444 3386 2628 3454
use cut_M2M3_1x2 
transform 1 0 1432 0 1 3328
box 1432 3328 1500 3512
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7850
box 2444 7850 2628 7918
use cut_M2M3_1x2 
transform 1 0 1244 0 1 7792
box 1244 7792 1312 7976
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7630
box 2444 7630 2628 7698
use cut_M2M3_1x2 
transform 1 0 1056 0 1 7572
box 1056 7572 1124 7756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8730
box 2444 8730 2628 8798
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8672
box 1056 8672 1124 8856
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8070
box 2444 8070 2628 8138
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8012
box 1056 8012 1124 8196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8510
box 2444 8510 2628 8578
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8452
box 1056 8452 1124 8636
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7630
box 2444 7630 2628 7698
use cut_M2M3_1x2 
transform 1 0 1056 0 1 7572
box 1056 7572 1124 7756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8730
box 2444 8730 2628 8798
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8672
box 1056 8672 1124 8856
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8070
box 2444 8070 2628 8138
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8012
box 1056 8012 1124 8196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8510
box 2444 8510 2628 8578
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8452
box 1056 8452 1124 8636
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7630
box 2444 7630 2628 7698
use cut_M2M3_1x2 
transform 1 0 1056 0 1 7572
box 1056 7572 1124 7756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8730
box 2444 8730 2628 8798
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8672
box 1056 8672 1124 8856
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8070
box 2444 8070 2628 8138
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8012
box 1056 8012 1124 8196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8510
box 2444 8510 2628 8578
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8452
box 1056 8452 1124 8636
use cut_M1M3_2x1 
transform 1 0 2444 0 1 7630
box 2444 7630 2628 7698
use cut_M2M3_1x2 
transform 1 0 1056 0 1 7572
box 1056 7572 1124 7756
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8730
box 2444 8730 2628 8798
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8672
box 1056 8672 1124 8856
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8070
box 2444 8070 2628 8138
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8012
box 1056 8012 1124 8196
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8510
box 2444 8510 2628 8578
use cut_M2M3_1x2 
transform 1 0 1056 0 1 8452
box 1056 8452 1124 8636
use cut_M1M3_2x1 
transform 1 0 2444 0 1 8290
box 2444 8290 2628 8358
use cut_M2M3_1x2 
transform 1 0 868 0 1 8232
box 868 8232 936 8416
use cut_M1M3_2x1 
transform 1 0 2444 0 1 3826
box 2444 3826 2628 3894
use cut_M2M3_1x2 
transform 1 0 680 0 1 3768
box 680 3768 748 3952
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4046
box 2444 4046 2628 4114
use cut_M2M3_1x2 
transform 1 0 492 0 1 3988
box 492 3988 560 4172
use cut_M1M3_2x1 
transform 1 0 2444 0 1 3606
box 2444 3606 2628 3674
use cut_M2M3_1x2 
transform 1 0 304 0 1 3548
box 304 3548 372 3732
use cut_M1M3_2x1 
transform 1 0 2444 0 1 4266
box 2444 4266 2628 4334
use cut_M2M3_1x2 
transform 1 0 116 0 1 4208
box 116 4208 184 4392
use cut_M1M2_1x2 
transform 1 0 2756 0 1 3108
box 2756 3108 2824 3292
use cut_M1M2_1x2 
transform 1 0 2756 0 1 3108
box 2756 3108 2824 3292
<< labels >>
flabel m1 s 2188 4596 2248 11904 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew
flabel m1 s 2000 132 2060 11904 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew
flabel m1 s 1812 9060 1872 11904 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew
flabel m1 s 1624 1620 1684 11904 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew
flabel m1 s 1436 3328 1496 11904 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew
flabel m1 s 1248 7792 1308 11904 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew
flabel m1 s 1060 7572 1120 11904 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew
flabel m1 s 872 8232 932 11904 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew
flabel m1 s 684 3768 744 11904 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew
flabel m1 s 496 3988 556 11904 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew
flabel m1 s 308 3548 368 11904 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew
flabel m1 s 120 4208 180 11904 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew
flabel m1 s 2756 0 11336 68 0 FreeSans 400 0 0 0 AVSS
port 13 nsew
flabel m3 s 2756 10416 2824 11964 0 FreeSans 400 0 0 0 CTOP
port 14 nsew
<< end >>
