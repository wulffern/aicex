magic
tech sky130A
magscale 1 2
timestamp 1660666507
<< checkpaint >>
rect 0 0 76 200
<< m2 >>
rect 0 0 76 200
<< m3 >>
rect 0 0 76 200
<< v2 >>
rect 6 12 70 188
<< labels >>
<< end >>
