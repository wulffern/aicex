magic
tech sky130A
magscale 1 2
timestamp 1660244192
<< checkpaint >>
rect -768 -768 3288 19424
<< locali >>
rect 2664 -384 2904 19040
rect -384 -384 2904 -144
rect -384 18800 2904 19040
rect -384 -384 -144 19040
rect 2664 -384 2904 19040
rect 3048 -768 3288 19424
rect -768 -768 3288 -528
rect -768 19184 3288 19424
rect -768 -768 -528 19424
rect 3048 -768 3288 19424
rect 432 850 600 910
rect 600 586 864 646
rect 600 586 660 910
rect 636 998 816 1058
rect 636 2698 864 2758
rect 432 1202 636 1262
rect 636 4458 864 4518
rect 432 2962 636 3022
rect 636 6218 864 6278
rect 432 4722 636 4782
rect 636 7978 864 8038
rect 432 6482 636 6542
rect 636 9738 864 9798
rect 432 8242 636 8302
rect 636 11498 864 11558
rect 432 10002 636 10062
rect 636 13258 864 13318
rect 432 11762 636 11822
rect 636 15018 864 15078
rect 432 13522 636 13582
rect 636 16778 864 16838
rect 432 15282 636 15342
rect 636 18538 864 18598
rect 432 17042 636 17102
rect 636 998 696 18598
rect 756 938 864 998
rect -108 352 108 17116
rect 756 938 972 998
rect 324 498 540 558
<< m3 >>
rect 748 -384 964 704
rect 1540 -768 1756 704
<< m1 >>
rect 864 762 1032 822
rect 864 1114 1032 1174
rect 864 2874 1032 2934
rect 864 4634 1032 4694
rect 864 6394 1032 6454
rect 864 8154 1032 8214
rect 864 9914 1032 9974
rect 864 11674 1032 11734
rect 864 13434 1032 13494
rect 864 15194 1032 15254
rect 864 16954 1032 17014
rect 856 352 1032 412
rect 1032 352 1092 17022
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV xa00
transform 1 0 0 0 1 0
box 0 0 2520 352
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa10
transform 1 0 0 0 1 352
box 0 352 2520 704
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa20
transform 1 0 0 0 1 704
box 0 704 1260 1056
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa30
transform 1 0 0 0 1 1056
box 0 1056 1260 2816
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa31
transform 1 0 0 0 1 2816
box 0 2816 1260 4576
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa32
transform 1 0 0 0 1 4576
box 0 4576 1260 6336
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa33
transform 1 0 0 0 1 6336
box 0 6336 1260 8096
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa34
transform 1 0 0 0 1 8096
box 0 8096 1260 9856
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa35
transform 1 0 0 0 1 9856
box 0 9856 1260 11616
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa36
transform 1 0 0 0 1 11616
box 0 11616 1260 13376
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa37
transform 1 0 0 0 1 13376
box 0 13376 1260 15136
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa38
transform 1 0 0 0 1 15136
box 0 15136 1260 16896
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa39
transform 1 0 0 0 1 16896
box 0 16896 1260 18656
use cut_M1M4_2x1 
transform 1 0 756 0 1 -384
box 756 -384 956 -308
use cut_M1M4_2x1 
transform 1 0 1548 0 1 -768
box 1548 -768 1748 -692
use cut_M1M2_2x1 
transform 1 0 788 0 1 762
box 788 762 972 830
use cut_M1M2_2x1 
transform 1 0 788 0 1 1114
box 788 1114 972 1182
use cut_M1M2_2x1 
transform 1 0 788 0 1 2874
box 788 2874 972 2942
use cut_M1M2_2x1 
transform 1 0 788 0 1 4634
box 788 4634 972 4702
use cut_M1M2_2x1 
transform 1 0 788 0 1 6394
box 788 6394 972 6462
use cut_M1M2_2x1 
transform 1 0 788 0 1 8154
box 788 8154 972 8222
use cut_M1M2_2x1 
transform 1 0 788 0 1 9914
box 788 9914 972 9982
use cut_M1M2_2x1 
transform 1 0 788 0 1 11674
box 788 11674 972 11742
use cut_M1M2_2x1 
transform 1 0 788 0 1 13434
box 788 13434 972 13502
use cut_M1M2_2x1 
transform 1 0 788 0 1 15194
box 788 15194 972 15262
use cut_M1M2_2x1 
transform 1 0 788 0 1 16954
box 788 16954 972 17022
use cut_M1M4_1x2 
transform 1 0 -38 0 1 352
box -38 352 38 552
<< labels >>
flabel locali s 2664 -384 2904 19040 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
flabel locali s 3048 -768 3288 19424 0 FreeSans 400 0 0 0 AVDD
port 2 nsew
flabel locali s 756 938 972 998 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
<< end >>
