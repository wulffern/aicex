magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 4480
<< locali >>
rect 1380 210 1534 270
rect 1534 710 1710 770
rect 1534 210 1594 770
rect 1650 770 1740 830
rect 1380 850 1534 910
rect 1534 1410 1740 1470
rect 1534 3970 1740 4030
rect 1534 850 1594 4030
rect 360 2050 514 2110
rect 514 850 720 910
rect 514 850 574 2110
rect 390 2950 514 3010
rect 514 850 720 910
rect 514 850 574 3010
rect 360 3010 450 3070
rect 720 1490 874 1550
rect 720 2130 874 2190
rect 874 1490 934 2190
rect 360 4290 514 4350
rect 514 4050 720 4110
rect 514 4050 574 4350
rect 270 1090 450 1150
rect 270 130 450 190
rect 630 4370 810 4430
rect 630 4050 810 4110
rect 270 3330 450 3390
rect 2010 120 2190 200
rect -90 120 90 200
<< m1 >>
rect 1740 2050 1894 2110
rect 1740 3010 1894 3070
rect 1380 210 1894 270
rect 1894 210 1954 3078
rect 390 1350 514 1410
rect 514 530 720 590
rect 514 530 574 1478
rect 360 1410 450 1470
rect 720 3090 874 3150
rect 720 4050 874 4110
rect 874 3090 934 4118
rect 360 2370 514 2430
rect 514 2130 720 2190
rect 514 2130 574 2438
rect 1380 2450 1534 2510
rect 1534 1730 1740 1790
rect 1534 2690 1740 2750
rect 1534 1730 1594 2758
rect 1380 4370 1534 4430
rect 1534 3650 1740 3710
rect 1534 3650 1594 4438
rect 146 450 360 510
rect 146 3330 360 3390
rect 146 450 206 3398
<< m2 >>
rect 360 3970 514 4038
rect 514 3010 1740 3078
rect 514 3010 582 4038
<< m3 >>
rect 1290 0 1474 4480
rect 630 0 814 4480
rect 1290 0 1474 4480
rect 630 0 814 4480
use NDX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2100 640
use IVX1_CV XA2
transform 1 0 0 0 1 640
box 0 640 2100 960
use IVTRIX1_CV XA3
transform 1 0 0 0 1 960
box 0 960 2100 1600
use IVTRIX1_CV XA4
transform 1 0 0 0 1 1600
box 0 1600 2100 2240
use IVX1_CV XA5
transform 1 0 0 0 1 2240
box 0 2240 2100 2560
use IVTRIX1_CV XA6
transform 1 0 0 0 1 2560
box 0 2560 2100 3200
use NDTRIX1_CV XA7
transform 1 0 0 0 1 3200
box 0 3200 2100 4160
use IVX1_CV XA8
transform 1 0 0 0 1 4160
box 0 4160 2100 4480
use cut_M1M2_2x1 
transform 1 0 1650 0 1 2050
box 1650 2050 1834 2118
use cut_M1M2_2x1 
transform 1 0 1650 0 1 3010
box 1650 3010 1834 3078
use cut_M1M2_2x1 
transform 1 0 1290 0 1 210
box 1290 210 1474 278
use cut_M1M2_2x1 
transform 1 0 270 0 1 1410
box 270 1410 454 1478
use cut_M1M2_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M3_2x1 
transform 1 0 270 0 1 3970
box 270 3970 454 4038
use cut_M1M3_2x1 
transform 1 0 1650 0 1 3010
box 1650 3010 1834 3078
use cut_M1M2_2x1 
transform 1 0 630 0 1 3090
box 630 3090 814 3158
use cut_M1M2_2x1 
transform 1 0 630 0 1 4050
box 630 4050 814 4118
use cut_M1M2_2x1 
transform 1 0 270 0 1 2370
box 270 2370 454 2438
use cut_M1M2_2x1 
transform 1 0 630 0 1 2130
box 630 2130 814 2198
use cut_M1M2_2x1 
transform 1 0 1290 0 1 2450
box 1290 2450 1474 2518
use cut_M1M2_2x1 
transform 1 0 1650 0 1 1730
box 1650 1730 1834 1798
use cut_M1M2_2x1 
transform 1 0 1650 0 1 2690
box 1650 2690 1834 2758
use cut_M1M2_2x1 
transform 1 0 1290 0 1 4370
box 1290 4370 1474 4438
use cut_M1M2_2x1 
transform 1 0 1650 0 1 3650
box 1650 3650 1834 3718
use cut_M1M2_2x1 
transform 1 0 270 0 1 450
box 270 450 454 518
use cut_M1M2_2x1 
transform 1 0 270 0 1 3330
box 270 3330 454 3398
<< labels >>
flabel locali s 270 1090 450 1150 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 CK
port 2 nsew
flabel locali s 630 4370 810 4430 0 FreeSans 400 0 0 0 Q
port 3 nsew
flabel locali s 630 4050 810 4110 0 FreeSans 400 0 0 0 QN
port 4 nsew
flabel locali s 270 3330 450 3390 0 FreeSans 400 0 0 0 RN
port 5 nsew
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 6 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 7 nsew
flabel m3 s 1290 0 1474 4480 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 4480 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
