magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect -5892 -2040 28148 39862
<< m3 >>
rect 8580 17864 26150 17924
rect 8580 18220 26150 18280
rect 22208 18552 22268 25432
rect 22496 18552 22556 32472
rect 3648 18636 3708 28628
rect 4488 18814 4548 28628
rect 8288 18992 8348 28628
rect -152 19170 -92 28628
rect 12324 19348 12384 28642
rect 16964 19526 17024 28642
rect 9864 19704 9924 28642
rect 14504 19882 14564 28642
rect 584 20060 644 28642
rect 5224 20238 5284 28642
rect 3044 20416 3104 28642
rect 7684 20594 7744 28642
rect 720 20772 780 29922
rect 7548 20950 7608 29922
rect 5360 21128 5420 29922
rect 2908 21306 2968 29922
rect 10136 21484 10196 31202
rect 12052 21662 12112 31202
rect 14776 21840 14836 31202
rect 7412 22018 7472 31202
rect 2772 22196 2832 31202
rect 856 22374 916 31202
rect 16692 22552 16752 31202
rect 5496 22730 5556 31202
rect 208 23382 408 38262
rect 3288 23382 3488 38262
rect 4848 23382 5048 38262
rect 7928 23382 8128 38262
rect 9488 23382 9688 38262
rect 12568 23382 12768 38262
rect 14128 23382 14328 38262
rect 17208 23382 17408 38262
rect 18768 23382 18968 38262
rect 21848 23382 22048 38262
rect 8888 -800 9088 4800
rect 13168 -800 13368 4800
rect 928 23382 1128 39062
rect 2568 23382 2768 39062
rect 5568 23382 5768 39062
rect 7208 23382 7408 39062
rect 10208 23382 10408 39062
rect 11848 23382 12048 39062
rect 14848 23382 15048 39062
rect 16488 23382 16688 39062
rect 19488 23382 19688 39062
rect 21128 23382 21328 39062
rect 8168 -1600 8368 4800
rect 13888 -1600 14088 4800
rect 1568 27752 1768 39862
rect 1928 27752 2128 39862
rect 6208 27752 6408 39862
rect 6568 27752 6768 39862
rect 10848 27752 11048 39862
rect 11208 27752 11408 39862
rect 15488 27752 15688 39862
rect 15848 27752 16048 39862
rect 20128 27752 20328 39862
rect 9518 -2040 9578 3154
rect 12678 -2040 12738 3154
rect 10100 1170 10328 1230
rect 8614 4978 10100 5038
rect 11928 1170 12096 1230
rect 12096 4978 13638 5038
rect 10328 1170 10496 1230
rect 10496 2450 11928 2510
rect 10496 1170 10556 2518
<< m2 >>
rect 13604 17390 13664 17932
rect 8580 17390 8640 18288
rect 3648 18576 12832 18636
rect 4488 18754 12520 18814
rect 8288 18932 12208 18992
rect -152 19110 13144 19170
rect 10512 19288 12384 19348
rect 10824 19466 17024 19526
rect 9864 19644 10416 19704
rect 10668 19822 14564 19882
rect 584 20000 9168 20060
rect 5224 20178 9792 20238
rect 3044 20356 9480 20416
rect 7684 20534 10104 20594
rect 720 20712 9324 20772
rect 7548 20890 10260 20950
rect 5360 21068 9948 21128
rect 2908 21246 9636 21306
rect 10136 21424 11896 21484
rect 11680 21602 12112 21662
rect 11524 21780 14836 21840
rect 7412 21958 12052 22018
rect 2772 22136 12676 22196
rect 856 22314 12988 22374
rect 11368 22492 16752 22552
rect 5496 22670 12364 22730
rect 928 36102 1264 36162
rect 1264 35564 3648 35624
rect 3588 35564 3648 35732
rect 1264 35564 1324 36174
rect 5568 36102 5904 36162
rect 5904 35564 8288 35624
rect 8228 35564 8288 35732
rect 5904 35564 5964 36174
rect 10208 36102 10544 36162
rect 10544 35564 12928 35624
rect 12868 35564 12928 35732
rect 10544 35564 10604 36174
rect 14848 36102 15184 36162
rect 15184 35564 17568 35624
rect 17508 35564 17568 35732
rect 15184 35564 15244 36174
rect -192 32684 18608 32744
rect -252 32684 -192 32852
rect 3588 32684 3648 32852
rect 4388 32684 4448 32852
rect 8228 32684 8288 32852
rect 9028 32684 9088 32852
rect 12868 32684 12928 32852
rect 13668 32684 13728 32852
rect 17508 32684 17568 32852
rect 18308 32684 18368 32852
rect 968 24068 1264 24128
rect 1264 23720 3648 23780
rect 3588 23720 3648 23896
rect 1264 23720 1324 24128
rect 5608 24068 5904 24128
rect 5904 23720 8288 23780
rect 8228 23720 8288 23896
rect 5904 23720 5964 24128
rect 10248 24068 10544 24128
rect 10544 23720 12928 23780
rect 12868 23720 12928 23896
rect 10544 23720 10604 24128
rect 14888 24068 15184 24128
rect 15184 23720 17568 23780
rect 17508 23720 17568 23896
rect 15184 23720 15244 24128
rect 19528 24068 19824 24128
rect 19824 24068 19884 24128
rect 2528 24068 2824 24128
rect 2824 24068 2884 24176
rect 2824 24176 4488 24236
rect 4428 23828 4488 24236
rect 7168 24068 7464 24128
rect 7464 24068 7524 24176
rect 7464 24176 9128 24236
rect 9068 23828 9128 24236
rect 11808 24068 12104 24128
rect 12104 24068 12164 24176
rect 12104 24176 13768 24236
rect 13708 23828 13768 24236
rect 16448 24068 16744 24128
rect 16744 24068 16804 24176
rect 16744 24176 18408 24236
rect 18348 23828 18408 24236
rect -152 25752 18608 25812
rect -212 25428 -152 25812
rect 3588 25428 3648 25812
rect 4428 25428 4488 25812
rect 8228 25428 8288 25812
rect 9068 25428 9128 25812
rect 12868 25428 12928 25812
rect 13708 25428 13768 25812
rect 17508 25428 17568 25812
rect 18348 25428 18408 25812
rect -192 26076 18608 26136
rect -252 26076 -192 26452
rect 3588 26076 3648 26452
rect 4388 26076 4448 26452
rect 8228 26076 8288 26452
rect 9028 26076 9088 26452
rect 12868 26076 12928 26452
rect 13668 26076 13728 26452
rect 17508 26076 17568 26452
rect 18308 26076 18368 26452
rect 1328 27032 48 27092
rect 1328 27032 1568 27092
rect 1328 27032 2368 27092
rect 1328 27032 6208 27092
rect 1328 27032 7008 27092
rect 1328 27032 10848 27092
rect 1328 27032 11648 27092
rect 1328 27032 15488 27092
rect 1328 27032 16288 27092
rect 1328 27032 20128 27092
rect 21700 28422 21928 28482
rect 18548 25488 21700 25548
rect 21700 25488 21760 28494
rect 18508 25428 18608 25488
rect 20980 29702 21208 29762
rect 18548 26452 20980 26512
rect 20980 26452 21040 29774
rect 18488 26392 18608 26452
rect 20808 36312 20976 36372
rect 18488 33432 20976 33492
rect 20976 33432 21036 36380
rect 20580 36952 20808 37012
rect 19608 36102 20580 36162
rect 20580 36102 20640 37020
rect 10328 2450 10496 2510
rect 10496 1170 11928 1230
rect 10496 1170 10556 2518
rect -192 27032 1568 27092
<< m4 >>
rect 22208 18220 22268 18552
rect 22496 17864 22556 18552
rect 10100 1170 10160 5038
rect 12096 1170 12156 5038
<< m1 >>
rect 12772 17330 12832 18576
rect 12460 17330 12520 18754
rect 12148 17330 12208 18932
rect 13084 17330 13144 19110
rect 10512 17330 10572 19288
rect 10824 17330 10884 19466
rect 10356 17330 10416 19644
rect 10668 17330 10728 19822
rect 9108 17330 9168 20000
rect 9732 17330 9792 20178
rect 9420 17330 9480 20356
rect 10044 17330 10104 20534
rect 9264 17330 9324 20712
rect 10200 17330 10260 20890
rect 9888 17330 9948 21068
rect 9576 17330 9636 21246
rect 11836 17330 11896 21424
rect 11680 17330 11740 21602
rect 11524 17330 11584 21780
rect 11992 17330 12052 21958
rect 12616 17330 12676 22136
rect 12928 17330 12988 22314
rect 11368 17330 11428 22492
rect 12304 17330 12364 22670
rect 9338 -1820 9398 510
rect 12858 -1820 12918 510
rect -192 35672 -5832 35732
rect 2528 36072 2864 36132
rect 2864 35564 4448 35624
rect 4388 35564 4448 35732
rect 2864 35564 2924 36140
rect 7168 36072 7504 36132
rect 7504 35564 9088 35624
rect 9028 35564 9088 35732
rect 7504 35564 7564 36140
rect 11808 36072 12144 36132
rect 12144 35564 13728 35624
rect 13668 35564 13728 35732
rect 12144 35564 12204 36140
rect 16448 36072 16784 36132
rect 16784 35564 18368 35624
rect 18308 35564 18368 35732
rect 16784 35564 16844 36140
rect 20580 36632 20808 36692
rect 18888 34152 20580 34212
rect 20580 34152 20640 36700
rect -4872 4978 68 5038
rect -4872 6522 68 6582
rect -4872 8066 68 8126
rect -4872 9610 68 9670
rect -4872 11154 68 11214
rect -4872 12698 68 12758
rect -4872 14242 68 14302
rect -4872 15786 68 15846
rect 22184 4978 27128 5038
rect 22184 6522 27128 6582
rect 22184 8066 27128 8126
rect 22184 9610 27128 9670
rect 22184 11154 27128 11214
rect 22184 12698 27128 12758
rect 22184 14242 27128 14302
rect 22184 15786 27128 15846
<< locali >>
rect -4872 -800 27128 -600
rect -4872 38062 27128 38262
rect -4872 -800 -4672 38262
rect 26928 -800 27128 38262
rect -5672 -1600 27928 -1400
rect -5672 38862 27928 39062
rect -5672 -1600 -5472 39062
rect 27728 -1600 27928 39062
rect -5672 39662 27928 39862
rect -5672 -1820 28148 -1760
rect 28088 -1820 28148 39862
rect -5892 -2040 28148 -1980
rect -5892 -2040 -5832 39862
use SARBSSW_CV XB1
transform -1 0 11128 0 1 0
box 11128 0 26328 4800
use SARBSSW_CV XB2
transform 1 0 11128 0 1 0
box 11128 0 26328 4800
use CDAC8_CV XDAC1
transform -1 0 11004 0 1 4978
box 11004 4978 21892 17390
use CDAC8_CV XDAC2
transform 1 0 11248 0 1 4978
box 11248 4978 22136 17390
use SARDIGEX4_CV XA0
transform 1 0 -472 0 1 23382
box -472 23382 1848 36502
use SARDIGEX4_CV XA1
transform -1 0 4168 0 1 23382
box 4168 23382 6488 36502
use SARDIGEX4_CV XA2
transform 1 0 4168 0 1 23382
box 4168 23382 6488 36502
use SARDIGEX4_CV XA3
transform -1 0 8808 0 1 23382
box 8808 23382 11128 36502
use SARDIGEX4_CV XA4
transform 1 0 8808 0 1 23382
box 8808 23382 11128 36502
use SARDIGEX4_CV XA5
transform -1 0 13448 0 1 23382
box 13448 23382 15768 36502
use SARDIGEX4_CV XA6
transform 1 0 13448 0 1 23382
box 13448 23382 15768 36502
use SARDIGEX4_CV XA7
transform -1 0 18088 0 1 23382
box 18088 23382 20408 36502
use SARDIGEX4_CV XA8
transform 1 0 18088 0 1 23382
box 18088 23382 20408 36502
use SARCMPX1_CV XA20
transform -1 0 22728 0 1 23382
box 22728 23382 25048 37462
use cut_M3M4_1x2 
transform 1 0 13604 0 1 17390
box 13604 17390 13672 17590
use cut_M3M4_2x1 
transform 1 0 13604 0 1 17864
box 13604 17864 13804 17932
use cut_M3M4_1x2 
transform 1 0 8580 0 1 17390
box 8580 17390 8648 17590
use cut_M3M4_2x1 
transform 1 0 8580 0 1 18220
box 8580 18220 8780 18288
use cut_M2M4_2x1 
transform 1 0 22208 0 1 25432
box 22208 25432 22408 25500
use cut_M4M5_2x1 
transform 1 0 22208 0 1 18220
box 22208 18220 22408 18288
use cut_M4M5_1x2 
transform 1 0 22208 0 1 18552
box 22208 18552 22276 18752
use cut_M3M4_2x1 
transform 1 0 22356 0 1 32472
box 22356 32472 22556 32540
use cut_M2M3_2x1 
transform 1 0 22208 0 1 32472
box 22208 32472 22408 32540
use cut_M4M5_2x1 
transform 1 0 22496 0 1 17864
box 22496 17864 22696 17932
use cut_M4M5_1x2 
transform 1 0 22496 0 1 18552
box 22496 18552 22564 18752
use cut_M3M4_1x2 
transform 1 0 3644 0 1 18506
box 3644 18506 3712 18706
use cut_M2M3_1x2 
transform 1 0 12768 0 1 18506
box 12768 18506 12836 18706
use cut_M3M4_1x2 
transform 1 0 4484 0 1 18684
box 4484 18684 4552 18884
use cut_M2M3_1x2 
transform 1 0 12456 0 1 18684
box 12456 18684 12524 18884
use cut_M3M4_1x2 
transform 1 0 8284 0 1 18862
box 8284 18862 8352 19062
use cut_M2M3_1x2 
transform 1 0 12144 0 1 18862
box 12144 18862 12212 19062
use cut_M3M4_1x2 
transform 1 0 -156 0 1 19040
box -156 19040 -88 19240
use cut_M2M3_1x2 
transform 1 0 13080 0 1 19040
box 13080 19040 13148 19240
use cut_M3M4_1x2 
transform 1 0 12320 0 1 19218
box 12320 19218 12388 19418
use cut_M2M3_1x2 
transform 1 0 10508 0 1 19218
box 10508 19218 10576 19418
use cut_M3M4_1x2 
transform 1 0 16960 0 1 19396
box 16960 19396 17028 19596
use cut_M2M3_1x2 
transform 1 0 10820 0 1 19396
box 10820 19396 10888 19596
use cut_M3M4_1x2 
transform 1 0 9860 0 1 19574
box 9860 19574 9928 19774
use cut_M2M3_1x2 
transform 1 0 10352 0 1 19574
box 10352 19574 10420 19774
use cut_M3M4_1x2 
transform 1 0 14500 0 1 19752
box 14500 19752 14568 19952
use cut_M2M3_1x2 
transform 1 0 10664 0 1 19752
box 10664 19752 10732 19952
use cut_M3M4_1x2 
transform 1 0 580 0 1 19930
box 580 19930 648 20130
use cut_M2M3_1x2 
transform 1 0 9104 0 1 19930
box 9104 19930 9172 20130
use cut_M3M4_1x2 
transform 1 0 5220 0 1 20108
box 5220 20108 5288 20308
use cut_M2M3_1x2 
transform 1 0 9728 0 1 20108
box 9728 20108 9796 20308
use cut_M3M4_1x2 
transform 1 0 3040 0 1 20286
box 3040 20286 3108 20486
use cut_M2M3_1x2 
transform 1 0 9416 0 1 20286
box 9416 20286 9484 20486
use cut_M3M4_1x2 
transform 1 0 7680 0 1 20464
box 7680 20464 7748 20664
use cut_M2M3_1x2 
transform 1 0 10040 0 1 20464
box 10040 20464 10108 20664
use cut_M3M4_1x2 
transform 1 0 716 0 1 20642
box 716 20642 784 20842
use cut_M2M3_1x2 
transform 1 0 9260 0 1 20642
box 9260 20642 9328 20842
use cut_M3M4_1x2 
transform 1 0 7544 0 1 20820
box 7544 20820 7612 21020
use cut_M2M3_1x2 
transform 1 0 10196 0 1 20820
box 10196 20820 10264 21020
use cut_M3M4_1x2 
transform 1 0 5356 0 1 20998
box 5356 20998 5424 21198
use cut_M2M3_1x2 
transform 1 0 9884 0 1 20998
box 9884 20998 9952 21198
use cut_M3M4_1x2 
transform 1 0 2904 0 1 21176
box 2904 21176 2972 21376
use cut_M2M3_1x2 
transform 1 0 9572 0 1 21176
box 9572 21176 9640 21376
use cut_M3M4_1x2 
transform 1 0 10132 0 1 21354
box 10132 21354 10200 21554
use cut_M2M3_1x2 
transform 1 0 11832 0 1 21354
box 11832 21354 11900 21554
use cut_M3M4_1x2 
transform 1 0 12048 0 1 21532
box 12048 21532 12116 21732
use cut_M2M3_1x2 
transform 1 0 11676 0 1 21532
box 11676 21532 11744 21732
use cut_M3M4_1x2 
transform 1 0 14772 0 1 21710
box 14772 21710 14840 21910
use cut_M2M3_1x2 
transform 1 0 11520 0 1 21710
box 11520 21710 11588 21910
use cut_M3M4_1x2 
transform 1 0 7408 0 1 21888
box 7408 21888 7476 22088
use cut_M2M3_1x2 
transform 1 0 11988 0 1 21888
box 11988 21888 12056 22088
use cut_M3M4_1x2 
transform 1 0 2768 0 1 22066
box 2768 22066 2836 22266
use cut_M2M3_1x2 
transform 1 0 12612 0 1 22066
box 12612 22066 12680 22266
use cut_M3M4_1x2 
transform 1 0 852 0 1 22244
box 852 22244 920 22444
use cut_M2M3_1x2 
transform 1 0 12924 0 1 22244
box 12924 22244 12992 22444
use cut_M3M4_1x2 
transform 1 0 16688 0 1 22422
box 16688 22422 16756 22622
use cut_M2M3_1x2 
transform 1 0 11364 0 1 22422
box 11364 22422 11432 22622
use cut_M3M4_1x2 
transform 1 0 5492 0 1 22600
box 5492 22600 5560 22800
use cut_M2M3_1x2 
transform 1 0 12300 0 1 22600
box 12300 22600 12368 22800
use cut_M1M4_2x2 
transform 1 0 208 0 1 38062
box 208 38062 408 38262
use cut_M1M4_2x2 
transform 1 0 3288 0 1 38062
box 3288 38062 3488 38262
use cut_M1M4_2x2 
transform 1 0 4848 0 1 38062
box 4848 38062 5048 38262
use cut_M1M4_2x2 
transform 1 0 7928 0 1 38062
box 7928 38062 8128 38262
use cut_M1M4_2x2 
transform 1 0 9488 0 1 38062
box 9488 38062 9688 38262
use cut_M1M4_2x2 
transform 1 0 12568 0 1 38062
box 12568 38062 12768 38262
use cut_M1M4_2x2 
transform 1 0 14128 0 1 38062
box 14128 38062 14328 38262
use cut_M1M4_2x2 
transform 1 0 17208 0 1 38062
box 17208 38062 17408 38262
use cut_M1M4_2x2 
transform 1 0 18768 0 1 38062
box 18768 38062 18968 38262
use cut_M1M4_2x2 
transform 1 0 21848 0 1 38062
box 21848 38062 22048 38262
use cut_M1M4_2x2 
transform 1 0 8888 0 1 -800
box 8888 -800 9088 -600
use cut_M1M4_2x2 
transform 1 0 13168 0 1 -800
box 13168 -800 13368 -600
use cut_M1M4_2x2 
transform 1 0 928 0 1 38862
box 928 38862 1128 39062
use cut_M1M4_2x2 
transform 1 0 2568 0 1 38862
box 2568 38862 2768 39062
use cut_M1M4_2x2 
transform 1 0 5568 0 1 38862
box 5568 38862 5768 39062
use cut_M1M4_2x2 
transform 1 0 7208 0 1 38862
box 7208 38862 7408 39062
use cut_M1M4_2x2 
transform 1 0 10208 0 1 38862
box 10208 38862 10408 39062
use cut_M1M4_2x2 
transform 1 0 11848 0 1 38862
box 11848 38862 12048 39062
use cut_M1M4_2x2 
transform 1 0 14848 0 1 38862
box 14848 38862 15048 39062
use cut_M1M4_2x2 
transform 1 0 16488 0 1 38862
box 16488 38862 16688 39062
use cut_M1M4_2x2 
transform 1 0 19488 0 1 38862
box 19488 38862 19688 39062
use cut_M1M4_2x2 
transform 1 0 21128 0 1 38862
box 21128 38862 21328 39062
use cut_M1M4_2x2 
transform 1 0 8168 0 1 -1600
box 8168 -1600 8368 -1400
use cut_M1M4_2x2 
transform 1 0 13888 0 1 -1600
box 13888 -1600 14088 -1400
use cut_M1M4_2x2 
transform 1 0 1568 0 1 39662
box 1568 39662 1768 39862
use cut_M1M4_2x2 
transform 1 0 1928 0 1 39662
box 1928 39662 2128 39862
use cut_M1M4_2x2 
transform 1 0 6208 0 1 39662
box 6208 39662 6408 39862
use cut_M1M4_2x2 
transform 1 0 6568 0 1 39662
box 6568 39662 6768 39862
use cut_M1M4_2x2 
transform 1 0 10848 0 1 39662
box 10848 39662 11048 39862
use cut_M1M4_2x2 
transform 1 0 11208 0 1 39662
box 11208 39662 11408 39862
use cut_M1M4_2x2 
transform 1 0 15488 0 1 39662
box 15488 39662 15688 39862
use cut_M1M4_2x2 
transform 1 0 15848 0 1 39662
box 15848 39662 16048 39862
use cut_M1M4_2x2 
transform 1 0 20128 0 1 39662
box 20128 39662 20328 39862
use cut_M1M2_2x1 
transform 1 0 9268 0 1 450
box 9268 450 9468 518
use cut_M1M2_2x1 
transform 1 0 9268 0 1 -1820
box 9268 -1820 9468 -1752
use cut_M1M2_2x1 
transform 1 0 12788 0 1 450
box 12788 450 12988 518
use cut_M1M2_2x1 
transform 1 0 12788 0 1 -1820
box 12788 -1820 12988 -1752
use cut_M1M2_2x1 
transform 1 0 -192 0 1 35672
box -192 35672 8 35740
use cut_M1M2_1x2 
transform 1 0 -5896 0 1 35602
box -5896 35602 -5828 35802
use cut_M1M4_2x1 
transform 1 0 9448 0 1 -2040
box 9448 -2040 9648 -1972
use cut_M1M4_2x1 
transform 1 0 12608 0 1 -2040
box 12608 -2040 12808 -1972
use cut_M1M3_2x1 
transform 1 0 928 0 1 36106
box 928 36106 1128 36174
use cut_M1M3_2x1 
transform 1 0 3648 0 1 35672
box 3648 35672 3848 35740
use cut_M1M3_2x1 
transform 1 0 5568 0 1 36106
box 5568 36106 5768 36174
use cut_M1M3_2x1 
transform 1 0 8288 0 1 35672
box 8288 35672 8488 35740
use cut_M1M3_2x1 
transform 1 0 10208 0 1 36106
box 10208 36106 10408 36174
use cut_M1M3_2x1 
transform 1 0 12928 0 1 35672
box 12928 35672 13128 35740
use cut_M1M3_2x1 
transform 1 0 14848 0 1 36106
box 14848 36106 15048 36174
use cut_M1M3_2x1 
transform 1 0 17568 0 1 35672
box 17568 35672 17768 35740
use cut_M1M3_2x1 
transform 1 0 -192 0 1 32792
box -192 32792 8 32860
use cut_M1M3_2x1 
transform 1 0 3648 0 1 32792
box 3648 32792 3848 32860
use cut_M1M3_2x1 
transform 1 0 4448 0 1 32792
box 4448 32792 4648 32860
use cut_M1M3_2x1 
transform 1 0 8288 0 1 32792
box 8288 32792 8488 32860
use cut_M1M3_2x1 
transform 1 0 9088 0 1 32792
box 9088 32792 9288 32860
use cut_M1M3_2x1 
transform 1 0 12928 0 1 32792
box 12928 32792 13128 32860
use cut_M1M3_2x1 
transform 1 0 13728 0 1 32792
box 13728 32792 13928 32860
use cut_M1M3_2x1 
transform 1 0 17568 0 1 32792
box 17568 32792 17768 32860
use cut_M1M3_2x1 
transform 1 0 18368 0 1 32792
box 18368 32792 18568 32860
use cut_M1M2_2x1 
transform 1 0 2528 0 1 36072
box 2528 36072 2728 36140
use cut_M1M2_2x1 
transform 1 0 4448 0 1 35672
box 4448 35672 4648 35740
use cut_M1M2_2x1 
transform 1 0 7168 0 1 36072
box 7168 36072 7368 36140
use cut_M1M2_2x1 
transform 1 0 9088 0 1 35672
box 9088 35672 9288 35740
use cut_M1M2_2x1 
transform 1 0 11808 0 1 36072
box 11808 36072 12008 36140
use cut_M1M2_2x1 
transform 1 0 13728 0 1 35672
box 13728 35672 13928 35740
use cut_M1M2_2x1 
transform 1 0 16448 0 1 36072
box 16448 36072 16648 36140
use cut_M1M2_2x1 
transform 1 0 18368 0 1 35672
box 18368 35672 18568 35740
use cut_M1M3_2x1 
transform 1 0 -192 0 1 26392
box -192 26392 8 26460
use cut_M1M3_2x1 
transform 1 0 3648 0 1 26392
box 3648 26392 3848 26460
use cut_M1M3_2x1 
transform 1 0 4448 0 1 26392
box 4448 26392 4648 26460
use cut_M1M3_2x1 
transform 1 0 8288 0 1 26392
box 8288 26392 8488 26460
use cut_M1M3_2x1 
transform 1 0 9088 0 1 26392
box 9088 26392 9288 26460
use cut_M1M3_2x1 
transform 1 0 12928 0 1 26392
box 12928 26392 13128 26460
use cut_M1M3_2x1 
transform 1 0 13728 0 1 26392
box 13728 26392 13928 26460
use cut_M1M3_2x1 
transform 1 0 17568 0 1 26392
box 17568 26392 17768 26460
use cut_M1M3_2x1 
transform 1 0 18368 0 1 26392
box 18368 26392 18568 26460
use cut_M1M3_2x1 
transform 1 0 1328 0 1 27032
box 1328 27032 1528 27100
use cut_M1M3_2x1 
transform 1 0 1328 0 1 27032
box 1328 27032 1528 27100
use cut_M1M3_2x1 
transform 1 0 2128 0 1 27032
box 2128 27032 2328 27100
use cut_M1M3_2x1 
transform 1 0 5968 0 1 27032
box 5968 27032 6168 27100
use cut_M1M3_2x1 
transform 1 0 6768 0 1 27032
box 6768 27032 6968 27100
use cut_M1M3_2x1 
transform 1 0 10608 0 1 27032
box 10608 27032 10808 27100
use cut_M1M3_2x1 
transform 1 0 11408 0 1 27032
box 11408 27032 11608 27100
use cut_M1M3_2x1 
transform 1 0 15248 0 1 27032
box 15248 27032 15448 27100
use cut_M1M3_2x1 
transform 1 0 16048 0 1 27032
box 16048 27032 16248 27100
use cut_M1M3_2x1 
transform 1 0 19888 0 1 27032
box 19888 27032 20088 27100
use cut_M1M3_2x1 
transform 1 0 21848 0 1 28426
box 21848 28426 22048 28494
use cut_M1M3_2x1 
transform 1 0 21128 0 1 29706
box 21128 29706 21328 29774
use cut_M1M3_2x1 
transform 1 0 20688 0 1 36312
box 20688 36312 20888 36380
use cut_M1M3_2x1 
transform 1 0 18368 0 1 33432
box 18368 33432 18568 33500
use cut_M1M3_2x1 
transform 1 0 20728 0 1 36952
box 20728 36952 20928 37020
use cut_M1M3_2x1 
transform 1 0 19528 0 1 36106
box 19528 36106 19728 36174
use cut_M1M2_2x1 
transform 1 0 20728 0 1 36632
box 20728 36632 20928 36700
use cut_M1M2_2x1 
transform 1 0 18808 0 1 34152
box 18808 34152 19008 34220
use cut_M4M5_1x2 
transform 1 0 10100 0 1 1170
box 10100 1170 10168 1370
use cut_M4M5_1x2 
transform 1 0 10100 0 1 4838
box 10100 4838 10168 5038
use cut_M1M4_2x1 
transform 1 0 11808 0 1 1170
box 11808 1170 12008 1238
use cut_M4M5_1x2 
transform 1 0 12096 0 1 1170
box 12096 1170 12164 1370
use cut_M4M5_1x2 
transform 1 0 12096 0 1 4838
box 12096 4838 12164 5038
use cut_M1M3_2x1 
transform 1 0 10208 0 1 2450
box 10208 2450 10408 2518
use cut_M1M3_2x1 
transform 1 0 11808 0 1 1170
box 11808 1170 12008 1238
use cut_M1M4_2x1 
transform 1 0 10208 0 1 1170
box 10208 1170 10408 1238
use cut_M1M4_2x1 
transform 1 0 11808 0 1 2450
box 11808 2450 12008 2518
use cut_M1M3_2x1 
transform 1 0 -192 0 1 27032
box -192 27032 8 27100
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 5038
box -4872 5038 -4672 5238
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 6582
box -4872 6582 -4672 6782
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 8126
box -4872 8126 -4672 8326
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 9670
box -4872 9670 -4672 9870
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 11214
box -4872 11214 -4672 11414
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 12758
box -4872 12758 -4672 12958
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 14302
box -4872 14302 -4672 14502
use cut_M1M2_2x2 
transform 1 0 -4872 0 1 15846
box -4872 15846 -4672 16046
use cut_M1M2_2x2 
transform 1 0 26928 0 1 4978
box 26928 4978 27128 5178
use cut_M1M2_2x2 
transform 1 0 26928 0 1 6522
box 26928 6522 27128 6722
use cut_M1M2_2x2 
transform 1 0 26928 0 1 8066
box 26928 8066 27128 8266
use cut_M1M2_2x2 
transform 1 0 26928 0 1 9610
box 26928 9610 27128 9810
use cut_M1M2_2x2 
transform 1 0 26928 0 1 11154
box 26928 11154 27128 11354
use cut_M1M2_2x2 
transform 1 0 26928 0 1 12698
box 26928 12698 27128 12898
use cut_M1M2_2x2 
transform 1 0 26928 0 1 14242
box 26928 14242 27128 14442
use cut_M1M2_2x2 
transform 1 0 26928 0 1 15786
box 26928 15786 27128 15986
<< labels >>
flabel m3 s -152 19170 -92 28628 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 12324 19348 12384 28642 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 16964 19526 17024 28642 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 9864 19704 9924 28642 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 14504 19882 14564 28642 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 5224 20238 5284 28642 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 3044 20416 3104 28642 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 7684 20594 7744 28642 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel locali s 26928 -800 27128 38262 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
flabel locali s 27728 -1600 27928 39062 0 FreeSans 400 0 0 0 AVDD
port 10 nsew
flabel locali s -5672 39662 27928 39862 0 FreeSans 400 0 0 0 VREF
port 11 nsew
flabel locali s 28088 -1820 28148 39862 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 12 nsew
flabel locali s 18768 34152 19008 34212 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 10208 46 10408 114 0 FreeSans 400 0 0 0 SAR_IP
port 14 nsew
flabel m3 s 11848 46 12048 114 0 FreeSans 400 0 0 0 SAR_IN
port 15 nsew
flabel locali s -192 32792 48 32852 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 1328 27032 1568 27092 0 FreeSans 400 0 0 0 EN
port 17 nsew
flabel locali s 10208 2450 10448 2510 0 FreeSans 400 0 0 0 SARN
port 18 nsew
flabel locali s 10208 1170 10448 1230 0 FreeSans 400 0 0 0 SARP
port 19 nsew
flabel m3 s 19144 28642 19212 28842 0 FreeSans 400 0 0 0 D<0>
port 20 nsew
<< end >>
