magic
tech sky130A
magscale 1 2
timestamp 1658582973
<< checkpaint >>
rect 0 0 2520 15488
<< locali >>
rect 1656 4986 1824 5046
rect 1824 9650 2088 9710
rect 1824 6834 2088 6894
rect 1824 4986 1884 9710
rect 204 2610 432 2670
rect 204 2962 432 3022
rect 204 8242 432 8302
rect 204 12818 432 12878
rect 204 2610 264 12878
rect 432 12818 600 12878
rect 600 13258 864 13318
rect 600 12818 660 13318
rect 636 14490 864 14550
rect 432 13522 636 13582
rect 636 13522 696 14550
rect 1656 15018 1824 15078
rect 1824 13874 2088 13934
rect 1824 13874 1884 15078
rect 636 4458 864 4518
rect 636 9738 864 9798
rect 636 4458 696 9798
rect 324 14226 540 14286
rect 324 14930 540 14990
rect 324 14578 540 14638
rect 756 6922 972 6982
rect 756 5514 972 5574
rect 324 2258 540 2318
rect 324 10002 540 10062
<< m1 >>
rect 1656 9562 1824 9622
rect 1824 4722 2088 4782
rect 1824 5426 2088 5486
rect 1824 4722 1884 9630
rect 432 2258 600 2318
rect 432 3314 600 3374
rect 600 2258 660 3382
rect 432 10002 600 10062
rect 432 11058 600 11118
rect 600 10002 660 11126
rect 204 498 432 558
rect 204 10706 432 10766
rect 204 13170 432 13230
rect 204 498 264 13238
rect 432 13170 600 13230
rect 600 13962 864 14022
rect 600 13170 660 14030
<< m3 >>
rect 1548 0 1748 15488
rect 756 0 956 15488
rect 1548 0 1748 15488
rect 756 0 956 15488
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use TAPCELLB_CV XA0
transform 1 0 0 0 1 0
box 0 0 2520 352
use SARKICKHX1_CV XA1
transform 1 0 0 0 1 352
box 0 352 2520 2816
use SARCMPHX1_CV XA2
transform 1 0 0 0 1 2816
box 0 2816 2520 5280
use IVX4_CV XA2a
transform 1 0 0 0 1 5280
box 0 5280 2520 6688
use IVX4_CV XA3a
transform 1 0 0 0 1 6688
box 0 6688 2520 8096
use SARCMPHX1_CV XA3
transform 1 0 0 0 1 8096
box 0 8096 2520 10560
use SARKICKHX1_CV XA4
transform 1 0 0 0 1 10560
box 0 10560 2520 13024
use IVX1_CV XA9
transform 1 0 0 0 1 13024
box 0 13024 2520 13376
use NDX1_CV XA10
transform 1 0 0 0 1 13376
box 0 13376 2520 14080
use NRX1_CV XA11
transform 1 0 0 0 1 14080
box 0 14080 2520 14784
use IVX1_CV XA12
transform 1 0 0 0 1 14784
box 0 14784 2520 15136
use TAPCELLB_CV XA13
transform 1 0 0 0 1 15136
box 0 15136 2520 15488
use DMY_CV XA14
transform 1 0 0 0 1 15488
box 0 15488 0 15488
use cut_M1M2_2x1 
transform 1 0 1548 0 1 9562
box 1548 9562 1732 9630
use cut_M1M2_2x1 
transform 1 0 1980 0 1 4722
box 1980 4722 2164 4790
use cut_M1M2_2x1 
transform 1 0 1980 0 1 5426
box 1980 5426 2164 5494
use cut_M1M2_2x1 
transform 1 0 356 0 1 2258
box 356 2258 540 2326
use cut_M1M2_2x1 
transform 1 0 356 0 1 3314
box 356 3314 540 3382
use cut_M1M2_2x1 
transform 1 0 356 0 1 10002
box 356 10002 540 10070
use cut_M1M2_2x1 
transform 1 0 356 0 1 11058
box 356 11058 540 11126
use cut_M1M2_2x1 
transform 1 0 324 0 1 498
box 324 498 508 566
use cut_M1M2_2x1 
transform 1 0 324 0 1 10706
box 324 10706 508 10774
use cut_M1M2_2x1 
transform 1 0 324 0 1 13170
box 324 13170 508 13238
use cut_M1M2_2x1 
transform 1 0 324 0 1 13170
box 324 13170 508 13238
use cut_M1M2_2x1 
transform 1 0 756 0 1 13962
box 756 13962 940 14030
<< labels >>
flabel locali s 324 14226 540 14286 0 FreeSans 400 0 0 0 CK_SAMPLE
port 1 nsew
flabel locali s 324 14930 540 14990 0 FreeSans 400 0 0 0 CK_CMP
port 2 nsew
flabel locali s 324 14578 540 14638 0 FreeSans 400 0 0 0 DONE
port 3 nsew
flabel locali s 756 6922 972 6982 0 FreeSans 400 0 0 0 CNO
port 4 nsew
flabel locali s 756 5514 972 5574 0 FreeSans 400 0 0 0 CPO
port 5 nsew
flabel locali s 324 2258 540 2318 0 FreeSans 400 0 0 0 CPI
port 6 nsew
flabel locali s 324 10002 540 10062 0 FreeSans 400 0 0 0 CNI
port 7 nsew
flabel m3 s 1548 0 1748 15488 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 756 0 956 15488 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
