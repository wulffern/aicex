magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect -3928 -1848 28016 57542
<< m3 >>
rect 9100 33880 26178 33956
rect 9100 34268 26178 34344
rect 24104 34648 24180 42152
rect 24384 34648 24460 49896
rect 3944 34732 4020 45664
rect 4824 34926 4900 45664
rect 8984 35120 9060 45664
rect -216 35314 -140 45664
rect -216 35314 -140 45664
rect 13432 35508 13508 45690
rect 13432 35508 13508 45690
rect 18472 35702 18548 45690
rect 18472 35702 18548 45690
rect 10579 35896 10655 45690
rect 10579 35896 10655 45690
rect 15619 36090 15695 45690
rect 15619 36090 15695 45690
rect 499 36284 575 45690
rect 5539 36478 5615 45690
rect 5539 36478 5615 45690
rect 3352 36672 3428 45690
rect 3352 36672 3428 45690
rect 8392 36866 8468 45690
rect 8392 36866 8468 45690
rect 659 37060 735 47098
rect 8232 37254 8308 47098
rect 5699 37448 5775 47098
rect 3192 37642 3268 47098
rect 10914 37836 10990 48506
rect 13098 38030 13174 48506
rect 15954 38224 16030 48506
rect 8058 38418 8134 48506
rect 3018 38612 3094 48506
rect 834 38806 910 48506
rect 18138 39000 18214 48506
rect 5874 39194 5950 48506
rect 200 39894 400 56102
rect 3528 39894 3728 56102
rect 5240 39894 5440 56102
rect 8568 39894 8768 56102
rect 10280 39894 10480 56102
rect 13608 39894 13808 56102
rect 15320 39894 15520 56102
rect 18648 39894 18848 56102
rect 20360 39894 20560 56102
rect 23688 39894 23888 56102
rect 9648 -720 9848 5280
rect 14240 -720 14440 5280
rect 992 39894 1192 56822
rect 2736 39894 2936 56822
rect 6032 39894 6232 56822
rect 7776 39894 7976 56822
rect 11072 39894 11272 56822
rect 12816 39894 13016 56822
rect 16112 39894 16312 56822
rect 17856 39894 18056 56822
rect 21152 39894 21352 56822
rect 22896 39894 23096 56822
rect 8856 -1440 9056 5280
rect 15032 -1440 15232 5280
rect 1568 44704 1768 57542
rect 2160 44704 2360 57542
rect 6608 44704 6808 57542
rect 7200 44704 7400 57542
rect 11648 44704 11848 57542
rect 12240 44704 12440 57542
rect 16688 44704 16888 57542
rect 17280 44704 17480 57542
rect 21728 44704 21928 57542
rect 10294 -1848 10370 3470
rect 13718 -1848 13794 3470
rect 10924 1290 11180 1366
rect 9138 5474 10924 5550
rect 12908 1290 13088 1366
rect 13088 5474 14910 5550
rect 11180 1290 11360 1366
rect 11360 2698 12908 2774
rect 11360 1290 11436 2774
rect 11072 50 11272 126
rect 12816 50 13016 126
rect 20659 45690 20735 45890
<< m2 >>
rect 14872 33374 14948 33956
rect 9100 33374 9176 34344
rect 3944 34656 14020 34732
rect 4824 34850 13660 34926
rect 8984 35044 13300 35120
rect -216 35238 14380 35314
rect 11304 35432 13508 35508
rect 11664 35626 18548 35702
rect 10579 35820 11200 35896
rect 11484 36014 15695 36090
rect 499 36208 9760 36284
rect 5539 36402 10480 36478
rect 3352 36596 10120 36672
rect 8392 36790 10840 36866
rect 659 36984 9940 37060
rect 8232 37178 11020 37254
rect 5699 37372 10660 37448
rect 3192 37566 10300 37642
rect 10914 37760 12940 37836
rect 12684 37954 13174 38030
rect 12504 38148 16030 38224
rect 8058 38342 13120 38418
rect 3018 38536 13840 38612
rect 834 38730 14200 38806
rect 12324 38924 18214 39000
rect 5874 39118 13480 39194
rect 992 53886 1336 53962
rect 1336 53276 3944 53352
rect 3868 53276 3944 53476
rect 1336 53276 1412 53970
rect 6032 53886 6376 53962
rect 6376 53276 8984 53352
rect 8908 53276 8984 53476
rect 6376 53276 6452 53970
rect 11072 53886 11416 53962
rect 11416 53276 14024 53352
rect 13948 53276 14024 53476
rect 11416 53276 11492 53970
rect 16112 53886 16456 53962
rect 16456 53276 19064 53352
rect 18988 53276 19064 53476
rect 16456 53276 16532 53970
rect -232 50108 20144 50184
rect -308 50108 -232 50308
rect 3868 50108 3944 50308
rect 4732 50108 4808 50308
rect 8908 50108 8984 50308
rect 9772 50108 9848 50308
rect 13948 50108 14024 50308
rect 14812 50108 14888 50308
rect 18988 50108 19064 50308
rect 19852 50108 19928 50308
rect 1008 40648 1336 40724
rect 1336 40244 3944 40320
rect 3868 40244 3944 40460
rect 1336 40244 1412 40724
rect 6048 40648 6376 40724
rect 6376 40244 8984 40320
rect 8908 40244 8984 40460
rect 6376 40244 6452 40724
rect 11088 40648 11416 40724
rect 11416 40244 14024 40320
rect 13948 40244 14024 40460
rect 11416 40244 11492 40724
rect 16128 40648 16456 40724
rect 16456 40244 19064 40320
rect 18988 40244 19064 40460
rect 16456 40244 16532 40724
rect 21168 40648 21496 40724
rect 21496 40648 21572 40724
rect 2720 40648 3048 40724
rect 3048 40648 3124 40788
rect 3048 40788 4824 40864
rect 4748 40384 4824 40864
rect 7760 40648 8088 40724
rect 8088 40648 8164 40788
rect 8088 40788 9864 40864
rect 9788 40384 9864 40864
rect 12800 40648 13128 40724
rect 13128 40648 13204 40788
rect 13128 40788 14904 40864
rect 14828 40384 14904 40864
rect 17840 40648 18168 40724
rect 18168 40648 18244 40788
rect 18168 40788 19944 40864
rect 19868 40384 19944 40864
rect -216 42436 20144 42512
rect -292 42144 -216 42512
rect 3868 42144 3944 42512
rect 4748 42144 4824 42512
rect 8908 42144 8984 42512
rect 9788 42144 9864 42512
rect 13948 42144 14024 42512
rect 14828 42144 14904 42512
rect 18988 42144 19064 42512
rect 19868 42144 19944 42512
rect -232 42916 20144 42992
rect -308 42916 -232 43268
rect 3868 42916 3944 43268
rect 4732 42916 4808 43268
rect 8908 42916 8984 43268
rect 9772 42916 9848 43268
rect 13948 42916 14024 43268
rect 14812 42916 14888 43268
rect 18988 42916 19064 43268
rect 19852 42916 19928 43268
rect -16 43912 1424 43972
rect 1424 43912 2504 43972
rect 1424 43912 6680 43972
rect 1424 43912 7544 43972
rect 1424 43912 11720 43972
rect 1424 43912 12584 43972
rect 1424 43912 16760 43972
rect 1424 43912 17624 43972
rect 1424 43912 21800 43972
rect 23396 45438 23780 45514
rect 20084 42220 23396 42296
rect 23396 42220 23472 45522
rect 20044 42144 20144 42220
rect 22740 46846 22988 46922
rect 20084 43284 22740 43360
rect 22740 43284 22816 46930
rect 20036 43208 20144 43284
rect 22556 54120 22728 54196
rect 20036 50952 22728 51028
rect 22728 50952 22804 54196
rect 22308 54824 22556 54900
rect 21260 53886 22308 53962
rect 22308 53886 22384 54900
rect 11180 2698 11352 2774
rect 11352 1290 12908 1366
rect 11352 1290 11428 2774
rect -232 43912 1640 43972
<< m4 >>
rect 24104 34268 24180 34648
rect 24384 33880 24460 34648
rect 10924 1290 11000 5550
rect 13088 1290 13164 5550
<< m1 >>
rect 13944 33314 14020 34656
rect 13584 33314 13660 34850
rect 13224 33314 13300 35044
rect 14304 33314 14380 35238
rect 11304 33314 11380 35432
rect 11664 33314 11740 35626
rect 11124 33314 11200 35820
rect 11484 33314 11560 36014
rect 9684 33314 9760 36208
rect 10404 33314 10480 36402
rect 10044 33314 10120 36596
rect 10764 33314 10840 36790
rect 9864 33314 9940 36984
rect 10944 33314 11020 37178
rect 10584 33314 10660 37372
rect 10224 33314 10300 37566
rect 12864 33314 12940 37760
rect 12684 33314 12760 37954
rect 12504 33314 12580 38148
rect 13044 33314 13120 38342
rect 13764 33314 13840 38536
rect 14124 33314 14200 38730
rect 12324 33314 12400 38924
rect 13404 33314 13480 39118
rect 10142 -1644 10202 558
rect 13886 -1644 13946 558
rect -3868 53416 -232 53476
rect 2720 53856 3056 53916
rect 3056 53296 4808 53356
rect 4748 53296 4808 53476
rect 3056 53296 3116 53924
rect 7760 53856 8096 53916
rect 8096 53296 9848 53356
rect 9788 53296 9848 53476
rect 8096 53296 8156 53924
rect 12800 53856 13136 53916
rect 13136 53296 14888 53356
rect 14828 53296 14888 53476
rect 13136 53296 13196 53924
rect 17840 53856 18176 53916
rect 18176 53296 19928 53356
rect 19868 53296 19928 53476
rect 18176 53296 18236 53924
rect 22328 54472 22556 54532
rect 20468 51744 22328 51804
rect 22328 51744 22388 54540
rect -3004 5474 76 5534
rect -3004 8954 76 9014
rect -3004 12434 76 12494
rect -3004 15914 76 15974
rect -3004 19394 76 19454
rect -3004 22874 76 22934
rect -3004 26354 76 26414
rect -3004 29834 76 29894
rect 23972 5474 27092 5534
rect 23972 8954 27092 9014
rect 23972 12434 27092 12494
rect 23972 15914 27092 15974
rect 23972 19394 27092 19454
rect 23972 22874 27092 22934
rect 23972 26354 27092 26414
rect 23972 29834 27092 29894
<< locali >>
rect 26892 -720 27092 56102
rect -3004 -720 27092 -520
rect -3004 55902 27092 56102
rect -3004 -720 -2804 56102
rect 26892 -720 27092 56102
rect 27612 -1440 27812 56822
rect -3724 -1440 27812 -1240
rect -3724 56622 27812 56822
rect -3724 -1440 -3524 56822
rect 27612 -1440 27812 56822
rect -3724 57342 27812 57542
rect -3724 57342 27812 57542
rect 27956 -1644 28016 57542
rect -3724 -1644 28016 -1584
rect 27956 -1644 28016 57542
rect -3928 -1848 28016 -1788
rect -3928 -1848 -3868 57542
rect 20360 51744 20576 51804
rect -232 50248 -16 50308
rect 1424 43912 1640 43972
rect 11072 2698 11288 2758
rect 11072 1290 11288 1350
use SUNSAR_SARBSSW_CV XB1
transform -1 0 12044 0 1 0
box 12044 0 26372 5280
use SUNSAR_SARBSSW_CV XB2
transform 1 0 12044 0 1 0
box 12044 0 26372 5280
use SUNSAR_CDAC8_CV XDAC1
transform -1 0 11844 0 1 5474
box 11844 5474 23576 33374
use SUNSAR_CDAC8_CV XDAC2
transform 1 0 12204 0 1 5474
box 12204 5474 23936 33374
use SUNSAR_SARDIGEX4_CV XA0
transform 1 0 -556 0 1 39894
box -556 39894 1964 54326
use SUNSAR_SARDIGEX4_CV XA1
transform -1 0 4484 0 1 39894
box 4484 39894 7004 54326
use SUNSAR_SARDIGEX4_CV XA2
transform 1 0 4484 0 1 39894
box 4484 39894 7004 54326
use SUNSAR_SARDIGEX4_CV XA3
transform -1 0 9524 0 1 39894
box 9524 39894 12044 54326
use SUNSAR_SARDIGEX4_CV XA4
transform 1 0 9524 0 1 39894
box 9524 39894 12044 54326
use SUNSAR_SARDIGEX4_CV XA5
transform -1 0 14564 0 1 39894
box 14564 39894 17084 54326
use SUNSAR_SARDIGEX4_CV XA6
transform 1 0 14564 0 1 39894
box 14564 39894 17084 54326
use SUNSAR_SARDIGEX4_CV XA7
transform -1 0 19604 0 1 39894
box 19604 39894 22124 54326
use SUNSAR_SARDIGEX4_CV XA8
transform 1 0 19604 0 1 39894
box 19604 39894 22124 54326
use SUNSAR_SARCMPX1_CV XA20
transform -1 0 24644 0 1 39894
box 24644 39894 27164 55382
use SUNSAR_cut_M3M4_1x2 
transform 1 0 14872 0 1 33374
box 14872 33374 14948 33574
use SUNSAR_cut_M3M4_2x1 
transform 1 0 14872 0 1 33880
box 14872 33880 15072 33956
use SUNSAR_cut_M3M4_1x2 
transform 1 0 9100 0 1 33374
box 9100 33374 9176 33574
use SUNSAR_cut_M3M4_2x1 
transform 1 0 9100 0 1 34268
box 9100 34268 9300 34344
use SUNSAR_cut_M2M4_2x1 
transform 1 0 24104 0 1 42152
box 24104 42152 24304 42228
use SUNSAR_cut_M4M5_2x1 
transform 1 0 24104 0 1 34268
box 24104 34268 24304 34344
use SUNSAR_cut_M4M5_1x2 
transform 1 0 24104 0 1 34648
box 24104 34648 24180 34848
use SUNSAR_cut_M3M4_2x1 
transform 1 0 24260 0 1 49896
box 24260 49896 24460 49972
use SUNSAR_cut_M2M3_2x1 
transform 1 0 24104 0 1 49896
box 24104 49896 24304 49972
use SUNSAR_cut_M4M5_2x1 
transform 1 0 24384 0 1 33880
box 24384 33880 24584 33956
use SUNSAR_cut_M4M5_1x2 
transform 1 0 24384 0 1 34648
box 24384 34648 24460 34848
use SUNSAR_cut_M3M4_1x2 
transform 1 0 3944 0 1 34594
box 3944 34594 4020 34794
use SUNSAR_cut_M2M3_1x2 
transform 1 0 13936 0 1 34594
box 13936 34594 14012 34794
use SUNSAR_cut_M3M4_1x2 
transform 1 0 4824 0 1 34788
box 4824 34788 4900 34988
use SUNSAR_cut_M2M3_1x2 
transform 1 0 13576 0 1 34788
box 13576 34788 13652 34988
use SUNSAR_cut_M3M4_1x2 
transform 1 0 8984 0 1 34982
box 8984 34982 9060 35182
use SUNSAR_cut_M2M3_1x2 
transform 1 0 13216 0 1 34982
box 13216 34982 13292 35182
use SUNSAR_cut_M3M4_1x2 
transform 1 0 -216 0 1 35176
box -216 35176 -140 35376
use SUNSAR_cut_M2M3_1x2 
transform 1 0 14296 0 1 35176
box 14296 35176 14372 35376
use SUNSAR_cut_M3M4_1x2 
transform 1 0 13432 0 1 35370
box 13432 35370 13508 35570
use SUNSAR_cut_M2M3_1x2 
transform 1 0 11296 0 1 35370
box 11296 35370 11372 35570
use SUNSAR_cut_M3M4_1x2 
transform 1 0 18472 0 1 35564
box 18472 35564 18548 35764
use SUNSAR_cut_M2M3_1x2 
transform 1 0 11656 0 1 35564
box 11656 35564 11732 35764
use SUNSAR_cut_M3M4_1x2 
transform 1 0 10579 0 1 35758
box 10579 35758 10655 35958
use SUNSAR_cut_M2M3_1x2 
transform 1 0 11116 0 1 35758
box 11116 35758 11192 35958
use SUNSAR_cut_M3M4_1x2 
transform 1 0 15619 0 1 35952
box 15619 35952 15695 36152
use SUNSAR_cut_M2M3_1x2 
transform 1 0 11476 0 1 35952
box 11476 35952 11552 36152
use SUNSAR_cut_M3M4_1x2 
transform 1 0 499 0 1 36146
box 499 36146 575 36346
use SUNSAR_cut_M2M3_1x2 
transform 1 0 9676 0 1 36146
box 9676 36146 9752 36346
use SUNSAR_cut_M3M4_1x2 
transform 1 0 5539 0 1 36340
box 5539 36340 5615 36540
use SUNSAR_cut_M2M3_1x2 
transform 1 0 10396 0 1 36340
box 10396 36340 10472 36540
use SUNSAR_cut_M3M4_1x2 
transform 1 0 3352 0 1 36534
box 3352 36534 3428 36734
use SUNSAR_cut_M2M3_1x2 
transform 1 0 10036 0 1 36534
box 10036 36534 10112 36734
use SUNSAR_cut_M3M4_1x2 
transform 1 0 8392 0 1 36728
box 8392 36728 8468 36928
use SUNSAR_cut_M2M3_1x2 
transform 1 0 10756 0 1 36728
box 10756 36728 10832 36928
use SUNSAR_cut_M3M4_1x2 
transform 1 0 659 0 1 36922
box 659 36922 735 37122
use SUNSAR_cut_M2M3_1x2 
transform 1 0 9856 0 1 36922
box 9856 36922 9932 37122
use SUNSAR_cut_M3M4_1x2 
transform 1 0 8232 0 1 37116
box 8232 37116 8308 37316
use SUNSAR_cut_M2M3_1x2 
transform 1 0 10936 0 1 37116
box 10936 37116 11012 37316
use SUNSAR_cut_M3M4_1x2 
transform 1 0 5699 0 1 37310
box 5699 37310 5775 37510
use SUNSAR_cut_M2M3_1x2 
transform 1 0 10576 0 1 37310
box 10576 37310 10652 37510
use SUNSAR_cut_M3M4_1x2 
transform 1 0 3192 0 1 37504
box 3192 37504 3268 37704
use SUNSAR_cut_M2M3_1x2 
transform 1 0 10216 0 1 37504
box 10216 37504 10292 37704
use SUNSAR_cut_M3M4_1x2 
transform 1 0 10914 0 1 37698
box 10914 37698 10990 37898
use SUNSAR_cut_M2M3_1x2 
transform 1 0 12856 0 1 37698
box 12856 37698 12932 37898
use SUNSAR_cut_M3M4_1x2 
transform 1 0 13098 0 1 37892
box 13098 37892 13174 38092
use SUNSAR_cut_M2M3_1x2 
transform 1 0 12676 0 1 37892
box 12676 37892 12752 38092
use SUNSAR_cut_M3M4_1x2 
transform 1 0 15954 0 1 38086
box 15954 38086 16030 38286
use SUNSAR_cut_M2M3_1x2 
transform 1 0 12496 0 1 38086
box 12496 38086 12572 38286
use SUNSAR_cut_M3M4_1x2 
transform 1 0 8058 0 1 38280
box 8058 38280 8134 38480
use SUNSAR_cut_M2M3_1x2 
transform 1 0 13036 0 1 38280
box 13036 38280 13112 38480
use SUNSAR_cut_M3M4_1x2 
transform 1 0 3018 0 1 38474
box 3018 38474 3094 38674
use SUNSAR_cut_M2M3_1x2 
transform 1 0 13756 0 1 38474
box 13756 38474 13832 38674
use SUNSAR_cut_M3M4_1x2 
transform 1 0 834 0 1 38668
box 834 38668 910 38868
use SUNSAR_cut_M2M3_1x2 
transform 1 0 14116 0 1 38668
box 14116 38668 14192 38868
use SUNSAR_cut_M3M4_1x2 
transform 1 0 18138 0 1 38862
box 18138 38862 18214 39062
use SUNSAR_cut_M2M3_1x2 
transform 1 0 12316 0 1 38862
box 12316 38862 12392 39062
use SUNSAR_cut_M3M4_1x2 
transform 1 0 5874 0 1 39056
box 5874 39056 5950 39256
use SUNSAR_cut_M2M3_1x2 
transform 1 0 13396 0 1 39056
box 13396 39056 13472 39256
use SUNSAR_cut_M1M4_2x2 
transform 1 0 200 0 1 55902
box 200 55902 400 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 3528 0 1 55902
box 3528 55902 3728 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 5240 0 1 55902
box 5240 55902 5440 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 8568 0 1 55902
box 8568 55902 8768 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 10280 0 1 55902
box 10280 55902 10480 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 13608 0 1 55902
box 13608 55902 13808 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 15320 0 1 55902
box 15320 55902 15520 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 18648 0 1 55902
box 18648 55902 18848 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 20360 0 1 55902
box 20360 55902 20560 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 23688 0 1 55902
box 23688 55902 23888 56102
use SUNSAR_cut_M1M4_2x2 
transform 1 0 9648 0 1 -720
box 9648 -720 9848 -520
use SUNSAR_cut_M1M4_2x2 
transform 1 0 14240 0 1 -720
box 14240 -720 14440 -520
use SUNSAR_cut_M1M4_2x2 
transform 1 0 992 0 1 56622
box 992 56622 1192 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 2736 0 1 56622
box 2736 56622 2936 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 6032 0 1 56622
box 6032 56622 6232 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 7776 0 1 56622
box 7776 56622 7976 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 11072 0 1 56622
box 11072 56622 11272 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 12816 0 1 56622
box 12816 56622 13016 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 16112 0 1 56622
box 16112 56622 16312 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 17856 0 1 56622
box 17856 56622 18056 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 21152 0 1 56622
box 21152 56622 21352 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 22896 0 1 56622
box 22896 56622 23096 56822
use SUNSAR_cut_M1M4_2x2 
transform 1 0 8856 0 1 -1440
box 8856 -1440 9056 -1240
use SUNSAR_cut_M1M4_2x2 
transform 1 0 15032 0 1 -1440
box 15032 -1440 15232 -1240
use SUNSAR_cut_M1M4_2x2 
transform 1 0 1568 0 1 57342
box 1568 57342 1768 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 2160 0 1 57342
box 2160 57342 2360 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 6608 0 1 57342
box 6608 57342 6808 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 7200 0 1 57342
box 7200 57342 7400 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 11648 0 1 57342
box 11648 57342 11848 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 12240 0 1 57342
box 12240 57342 12440 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 16688 0 1 57342
box 16688 57342 16888 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 17280 0 1 57342
box 17280 57342 17480 57542
use SUNSAR_cut_M1M4_2x2 
transform 1 0 21728 0 1 57342
box 21728 57342 21928 57542
use SUNSAR_cut_M1M2_2x1 
transform 1 0 10080 0 1 498
box 10080 498 10264 566
use SUNSAR_cut_M1M2_2x1 
transform 1 0 10080 0 1 -1644
box 10080 -1644 10264 -1576
use SUNSAR_cut_M1M2_2x1 
transform 1 0 13824 0 1 498
box 13824 498 14008 566
use SUNSAR_cut_M1M2_2x1 
transform 1 0 13824 0 1 -1644
box 13824 -1644 14008 -1576
use SUNSAR_cut_M1M2_2x1 
transform 1 0 -232 0 1 53416
box -232 53416 -48 53484
use SUNSAR_cut_M1M2_1x2 
transform 1 0 -3932 0 1 53354
box -3932 53354 -3864 53538
use SUNSAR_cut_M1M4_2x1 
transform 1 0 10232 0 1 -1848
box 10232 -1848 10432 -1772
use SUNSAR_cut_M1M4_2x1 
transform 1 0 13656 0 1 -1848
box 13656 -1848 13856 -1772
use SUNSAR_cut_M1M3_2x1 
transform 1 0 992 0 1 53894
box 992 53894 1192 53970
use SUNSAR_cut_M1M3_2x1 
transform 1 0 3944 0 1 53416
box 3944 53416 4144 53492
use SUNSAR_cut_M1M3_2x1 
transform 1 0 6032 0 1 53894
box 6032 53894 6232 53970
use SUNSAR_cut_M1M3_2x1 
transform 1 0 8984 0 1 53416
box 8984 53416 9184 53492
use SUNSAR_cut_M1M3_2x1 
transform 1 0 11072 0 1 53894
box 11072 53894 11272 53970
use SUNSAR_cut_M1M3_2x1 
transform 1 0 14024 0 1 53416
box 14024 53416 14224 53492
use SUNSAR_cut_M1M3_2x1 
transform 1 0 16112 0 1 53894
box 16112 53894 16312 53970
use SUNSAR_cut_M1M3_2x1 
transform 1 0 19064 0 1 53416
box 19064 53416 19264 53492
use SUNSAR_cut_M1M3_2x1 
transform 1 0 -232 0 1 50248
box -232 50248 -32 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 3944 0 1 50248
box 3944 50248 4144 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 4808 0 1 50248
box 4808 50248 5008 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 8984 0 1 50248
box 8984 50248 9184 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 9848 0 1 50248
box 9848 50248 10048 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 14024 0 1 50248
box 14024 50248 14224 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 14888 0 1 50248
box 14888 50248 15088 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 19064 0 1 50248
box 19064 50248 19264 50324
use SUNSAR_cut_M1M3_2x1 
transform 1 0 19928 0 1 50248
box 19928 50248 20128 50324
use SUNSAR_cut_M1M2_2x1 
transform 1 0 2720 0 1 53856
box 2720 53856 2904 53924
use SUNSAR_cut_M1M2_2x1 
transform 1 0 4808 0 1 53416
box 4808 53416 4992 53484
use SUNSAR_cut_M1M2_2x1 
transform 1 0 7760 0 1 53856
box 7760 53856 7944 53924
use SUNSAR_cut_M1M2_2x1 
transform 1 0 9848 0 1 53416
box 9848 53416 10032 53484
use SUNSAR_cut_M1M2_2x1 
transform 1 0 12800 0 1 53856
box 12800 53856 12984 53924
use SUNSAR_cut_M1M2_2x1 
transform 1 0 14888 0 1 53416
box 14888 53416 15072 53484
use SUNSAR_cut_M1M2_2x1 
transform 1 0 17840 0 1 53856
box 17840 53856 18024 53924
use SUNSAR_cut_M1M2_2x1 
transform 1 0 19928 0 1 53416
box 19928 53416 20112 53484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 -232 0 1 43208
box -232 43208 -32 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 3944 0 1 43208
box 3944 43208 4144 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 4808 0 1 43208
box 4808 43208 5008 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 8984 0 1 43208
box 8984 43208 9184 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 9848 0 1 43208
box 9848 43208 10048 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 14024 0 1 43208
box 14024 43208 14224 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 14888 0 1 43208
box 14888 43208 15088 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 19064 0 1 43208
box 19064 43208 19264 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 19928 0 1 43208
box 19928 43208 20128 43284
use SUNSAR_cut_M1M3_2x1 
transform 1 0 1424 0 1 43912
box 1424 43912 1624 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2288 0 1 43912
box 2288 43912 2488 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 6464 0 1 43912
box 6464 43912 6664 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 7328 0 1 43912
box 7328 43912 7528 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 11504 0 1 43912
box 11504 43912 11704 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 12368 0 1 43912
box 12368 43912 12568 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 16544 0 1 43912
box 16544 43912 16744 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 17408 0 1 43912
box 17408 43912 17608 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 21584 0 1 43912
box 21584 43912 21784 43988
use SUNSAR_cut_M1M3_2x1 
transform 1 0 23688 0 1 45446
box 23688 45446 23888 45522
use SUNSAR_cut_M1M3_2x1 
transform 1 0 22896 0 1 46854
box 22896 46854 23096 46930
use SUNSAR_cut_M1M3_2x1 
transform 1 0 22448 0 1 54120
box 22448 54120 22648 54196
use SUNSAR_cut_M1M3_2x1 
transform 1 0 19928 0 1 50952
box 19928 50952 20128 51028
use SUNSAR_cut_M1M3_2x1 
transform 1 0 22464 0 1 54824
box 22464 54824 22664 54900
use SUNSAR_cut_M1M3_2x1 
transform 1 0 21168 0 1 53894
box 21168 53894 21368 53970
use SUNSAR_cut_M1M2_2x1 
transform 1 0 22480 0 1 54472
box 22480 54472 22664 54540
use SUNSAR_cut_M1M2_2x1 
transform 1 0 20392 0 1 51744
box 20392 51744 20576 51812
use SUNSAR_cut_M4M5_1x2 
transform 1 0 10924 0 1 1290
box 10924 1290 11000 1490
use SUNSAR_cut_M4M5_1x2 
transform 1 0 10924 0 1 5350
box 10924 5350 11000 5550
use SUNSAR_cut_M1M4_2x1 
transform 1 0 12800 0 1 1290
box 12800 1290 13000 1366
use SUNSAR_cut_M4M5_1x2 
transform 1 0 13088 0 1 1290
box 13088 1290 13164 1490
use SUNSAR_cut_M4M5_1x2 
transform 1 0 13088 0 1 5350
box 13088 5350 13164 5550
use SUNSAR_cut_M1M3_2x1 
transform 1 0 11072 0 1 2698
box 11072 2698 11272 2774
use SUNSAR_cut_M1M3_2x1 
transform 1 0 12800 0 1 1290
box 12800 1290 13000 1366
use SUNSAR_cut_M1M4_2x1 
transform 1 0 11072 0 1 1290
box 11072 1290 11272 1366
use SUNSAR_cut_M1M4_2x1 
transform 1 0 12800 0 1 2698
box 12800 2698 13000 2774
use SUNSAR_cut_M1M3_2x1 
transform 1 0 -232 0 1 43912
box -232 43912 -32 43988
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 5534
box -3004 5534 -2820 5718
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 9014
box -3004 9014 -2820 9198
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 12494
box -3004 12494 -2820 12678
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 15974
box -3004 15974 -2820 16158
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 19454
box -3004 19454 -2820 19638
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 22934
box -3004 22934 -2820 23118
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 26414
box -3004 26414 -2820 26598
use SUNSAR_cut_M1M2_2x2 
transform 1 0 -3004 0 1 29894
box -3004 29894 -2820 30078
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 5474
box 27024 5474 27092 5658
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 8954
box 27024 8954 27092 9138
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 12434
box 27024 12434 27092 12618
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 15914
box 27024 15914 27092 16098
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 19394
box 27024 19394 27092 19578
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 22874
box 27024 22874 27092 23058
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 26354
box 27024 26354 27092 26538
use SUNSAR_cut_M1M2_1x2 
transform 1 0 27024 0 1 29834
box 27024 29834 27092 30018
<< labels >>
flabel m3 s -216 35314 -140 45664 0 FreeSans 400 0 0 0 D<8>
port 6 nsew
flabel m3 s 13432 35508 13508 45690 0 FreeSans 400 0 0 0 D<3>
port 11 nsew
flabel m3 s 18472 35702 18548 45690 0 FreeSans 400 0 0 0 D<1>
port 13 nsew
flabel m3 s 10579 35896 10655 45690 0 FreeSans 400 0 0 0 D<4>
port 10 nsew
flabel m3 s 15619 36090 15695 45690 0 FreeSans 400 0 0 0 D<2>
port 12 nsew
flabel m3 s 5539 36478 5615 45690 0 FreeSans 400 0 0 0 D<6>
port 8 nsew
flabel m3 s 3352 36672 3428 45690 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8392 36866 8468 45690 0 FreeSans 400 0 0 0 D<5>
port 9 nsew
flabel locali s 26892 -720 27092 56102 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
flabel locali s 27612 -1440 27812 56822 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel locali s -3724 57342 27812 57542 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel locali s 27956 -1644 28016 57542 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel locali s 20360 51744 20576 51804 0 FreeSans 400 0 0 0 DONE
port 5 nsew
flabel m3 s 11072 50 11272 126 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew
flabel m3 s 12816 50 13016 126 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew
flabel locali s -232 50248 -16 50308 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 1424 43912 1640 43972 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s 11072 2698 11288 2758 0 FreeSans 400 0 0 0 SARN
port 3 nsew
flabel locali s 11072 1290 11288 1350 0 FreeSans 400 0 0 0 SARP
port 4 nsew
flabel m3 s 20659 45690 20735 45890 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
<< end >>
