magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 116 0 11004 12412
<< m1 >>
rect 1836 4764 1896 12352
rect 1680 132 1740 12352
rect 1524 9396 1584 12352
rect 1368 1676 1428 12352
rect 1212 3448 1272 12352
rect 1056 8080 1116 12352
rect 900 7852 960 12352
rect 744 8536 804 12352
rect 588 3904 648 12352
rect 432 4132 492 12352
rect 276 3676 336 12352
rect 120 4360 180 12352
<< m2 >>
rect 2028 4830 1896 4898
rect 2028 5970 1896 6038
rect 2028 5286 1896 5354
rect 2028 5742 1896 5810
rect 2028 5514 1896 5582
rect 2028 5058 1896 5126
rect 2028 4830 1896 4898
rect 2028 5970 1896 6038
rect 2028 5286 1896 5354
rect 2028 5742 1896 5810
rect 2028 5514 1896 5582
rect 2028 5058 1896 5126
rect 2028 4830 1896 4898
rect 2028 5970 1896 6038
rect 2028 5286 1896 5354
rect 2028 5742 1896 5810
rect 2028 5514 1896 5582
rect 2028 5058 1896 5126
rect 2028 4830 1896 4898
rect 2028 5970 1896 6038
rect 2028 5286 1896 5354
rect 2028 5742 1896 5810
rect 2028 5514 1896 5582
rect 2028 5058 1896 5126
rect 2028 4830 1896 4898
rect 2028 5970 1896 6038
rect 2028 5286 1896 5354
rect 2028 5742 1896 5810
rect 2028 5514 1896 5582
rect 2028 5058 1896 5126
rect 2028 4830 1896 4898
rect 2028 5970 1896 6038
rect 2028 5286 1896 5354
rect 2028 5742 1896 5810
rect 2028 5514 1896 5582
rect 2028 5058 1896 5126
rect 2028 11006 1896 11074
rect 2028 12146 1896 12214
rect 2028 11462 1896 11530
rect 2028 11918 1896 11986
rect 2028 11690 1896 11758
rect 2028 11234 1896 11302
rect 2028 11006 1896 11074
rect 2028 12146 1896 12214
rect 2028 11462 1896 11530
rect 2028 11918 1896 11986
rect 2028 11690 1896 11758
rect 2028 11234 1896 11302
rect 2028 11006 1896 11074
rect 2028 12146 1896 12214
rect 2028 11462 1896 11530
rect 2028 11918 1896 11986
rect 2028 11690 1896 11758
rect 2028 11234 1896 11302
rect 2028 11006 1896 11074
rect 2028 12146 1896 12214
rect 2028 11462 1896 11530
rect 2028 11918 1896 11986
rect 2028 11690 1896 11758
rect 2028 11234 1896 11302
rect 2028 11006 1896 11074
rect 2028 12146 1896 12214
rect 2028 11462 1896 11530
rect 2028 11918 1896 11986
rect 2028 11690 1896 11758
rect 2028 11234 1896 11302
rect 2028 11006 1896 11074
rect 2028 12146 1896 12214
rect 2028 11462 1896 11530
rect 2028 11918 1896 11986
rect 2028 11690 1896 11758
rect 2028 11234 1896 11302
rect 2028 198 1740 266
rect 2028 1338 1740 1406
rect 2028 654 1740 722
rect 2028 1110 1740 1178
rect 2028 882 1740 950
rect 2028 426 1740 494
rect 2028 198 1740 266
rect 2028 1338 1740 1406
rect 2028 654 1740 722
rect 2028 1110 1740 1178
rect 2028 882 1740 950
rect 2028 426 1740 494
rect 2028 198 1740 266
rect 2028 1338 1740 1406
rect 2028 654 1740 722
rect 2028 1110 1740 1178
rect 2028 882 1740 950
rect 2028 426 1740 494
rect 2028 198 1740 266
rect 2028 1338 1740 1406
rect 2028 654 1740 722
rect 2028 1110 1740 1178
rect 2028 882 1740 950
rect 2028 426 1740 494
rect 2028 198 1740 266
rect 2028 1338 1740 1406
rect 2028 654 1740 722
rect 2028 1110 1740 1178
rect 2028 882 1740 950
rect 2028 426 1740 494
rect 2028 198 1740 266
rect 2028 1338 1740 1406
rect 2028 654 1740 722
rect 2028 1110 1740 1178
rect 2028 882 1740 950
rect 2028 426 1740 494
rect 2028 6374 1740 6442
rect 2028 7514 1740 7582
rect 2028 6830 1740 6898
rect 2028 7286 1740 7354
rect 2028 7058 1740 7126
rect 2028 6602 1740 6670
rect 2028 6374 1740 6442
rect 2028 7514 1740 7582
rect 2028 6830 1740 6898
rect 2028 7286 1740 7354
rect 2028 7058 1740 7126
rect 2028 6602 1740 6670
rect 2028 6374 1740 6442
rect 2028 7514 1740 7582
rect 2028 6830 1740 6898
rect 2028 7286 1740 7354
rect 2028 7058 1740 7126
rect 2028 6602 1740 6670
rect 2028 6374 1740 6442
rect 2028 7514 1740 7582
rect 2028 6830 1740 6898
rect 2028 7286 1740 7354
rect 2028 7058 1740 7126
rect 2028 6602 1740 6670
rect 2028 6374 1740 6442
rect 2028 7514 1740 7582
rect 2028 6830 1740 6898
rect 2028 7286 1740 7354
rect 2028 7058 1740 7126
rect 2028 6602 1740 6670
rect 2028 6374 1740 6442
rect 2028 7514 1740 7582
rect 2028 6830 1740 6898
rect 2028 7286 1740 7354
rect 2028 7058 1740 7126
rect 2028 6602 1740 6670
rect 2028 9462 1584 9530
rect 2028 10602 1584 10670
rect 2028 9918 1584 9986
rect 2028 10374 1584 10442
rect 2028 10146 1584 10214
rect 2028 9690 1584 9758
rect 2028 9462 1584 9530
rect 2028 10602 1584 10670
rect 2028 9918 1584 9986
rect 2028 10374 1584 10442
rect 2028 10146 1584 10214
rect 2028 9690 1584 9758
rect 2028 9462 1584 9530
rect 2028 10602 1584 10670
rect 2028 9918 1584 9986
rect 2028 10374 1584 10442
rect 2028 10146 1584 10214
rect 2028 9690 1584 9758
rect 2028 9462 1584 9530
rect 2028 10602 1584 10670
rect 2028 9918 1584 9986
rect 2028 10374 1584 10442
rect 2028 10146 1584 10214
rect 2028 9690 1584 9758
rect 2028 9462 1584 9530
rect 2028 10602 1584 10670
rect 2028 9918 1584 9986
rect 2028 10374 1584 10442
rect 2028 10146 1584 10214
rect 2028 9690 1584 9758
rect 2028 9462 1584 9530
rect 2028 10602 1584 10670
rect 2028 9918 1584 9986
rect 2028 10374 1584 10442
rect 2028 10146 1584 10214
rect 2028 9690 1584 9758
rect 2028 1742 1428 1810
rect 2028 2882 1428 2950
rect 2028 2198 1428 2266
rect 2028 2654 1428 2722
rect 2028 2426 1428 2494
rect 2028 1970 1428 2038
rect 2028 1742 1428 1810
rect 2028 2882 1428 2950
rect 2028 2198 1428 2266
rect 2028 2654 1428 2722
rect 2028 2426 1428 2494
rect 2028 1970 1428 2038
rect 2028 1742 1428 1810
rect 2028 2882 1428 2950
rect 2028 2198 1428 2266
rect 2028 2654 1428 2722
rect 2028 2426 1428 2494
rect 2028 1970 1428 2038
rect 2028 1742 1428 1810
rect 2028 2882 1428 2950
rect 2028 2198 1428 2266
rect 2028 2654 1428 2722
rect 2028 2426 1428 2494
rect 2028 1970 1428 2038
rect 2028 1742 1428 1810
rect 2028 2882 1428 2950
rect 2028 2198 1428 2266
rect 2028 2654 1428 2722
rect 2028 2426 1428 2494
rect 2028 1970 1428 2038
rect 2028 1742 1428 1810
rect 2028 2882 1428 2950
rect 2028 2198 1428 2266
rect 2028 2654 1428 2722
rect 2028 2426 1428 2494
rect 2028 1970 1428 2038
rect 2028 3514 1272 3582
rect 2028 8146 1116 8214
rect 2028 7918 960 7986
rect 2028 9058 960 9126
rect 2028 8374 960 8442
rect 2028 8830 960 8898
rect 2028 7918 960 7986
rect 2028 9058 960 9126
rect 2028 8374 960 8442
rect 2028 8830 960 8898
rect 2028 7918 960 7986
rect 2028 9058 960 9126
rect 2028 8374 960 8442
rect 2028 8830 960 8898
rect 2028 7918 960 7986
rect 2028 9058 960 9126
rect 2028 8374 960 8442
rect 2028 8830 960 8898
rect 2028 8602 804 8670
rect 2028 3970 648 4038
rect 2028 4198 492 4266
rect 2028 3742 336 3810
rect 2028 4426 180 4494
use CAP32C_CV XC1
transform 1 0 2028 0 1 0
box 2028 0 11004 1544
use CAP32C_CV XC64a<0>
transform 1 0 2028 0 1 1544
box 2028 1544 11004 3088
use CAP32C_CV XC32a<0>
transform 1 0 2028 0 1 3088
box 2028 3088 11004 4632
use CAP32C_CV XC128a<1>
transform 1 0 2028 0 1 4632
box 2028 4632 11004 6176
use CAP32C_CV XC128b<2>
transform 1 0 2028 0 1 6176
box 2028 6176 11004 7720
use CAP32C_CV X16ab
transform 1 0 2028 0 1 7720
box 2028 7720 11004 9264
use CAP32C_CV XC64b<1>
transform 1 0 2028 0 1 9264
box 2028 9264 11004 10808
use CAP32C_CV XC0
transform 1 0 2028 0 1 10808
box 2028 10808 11004 12352
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4830
box 2028 4830 2228 4898
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4764
box 1832 4764 1900 4964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5970
box 2028 5970 2228 6038
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5904
box 1832 5904 1900 6104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5286
box 2028 5286 2228 5354
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5220
box 1832 5220 1900 5420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5742
box 2028 5742 2228 5810
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5676
box 1832 5676 1900 5876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5514
box 2028 5514 2228 5582
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5448
box 1832 5448 1900 5648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5058
box 2028 5058 2228 5126
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4992
box 1832 4992 1900 5192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4830
box 2028 4830 2228 4898
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4764
box 1832 4764 1900 4964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5970
box 2028 5970 2228 6038
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5904
box 1832 5904 1900 6104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5286
box 2028 5286 2228 5354
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5220
box 1832 5220 1900 5420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5742
box 2028 5742 2228 5810
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5676
box 1832 5676 1900 5876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5514
box 2028 5514 2228 5582
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5448
box 1832 5448 1900 5648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5058
box 2028 5058 2228 5126
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4992
box 1832 4992 1900 5192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4830
box 2028 4830 2228 4898
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4764
box 1832 4764 1900 4964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5970
box 2028 5970 2228 6038
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5904
box 1832 5904 1900 6104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5286
box 2028 5286 2228 5354
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5220
box 1832 5220 1900 5420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5742
box 2028 5742 2228 5810
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5676
box 1832 5676 1900 5876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5514
box 2028 5514 2228 5582
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5448
box 1832 5448 1900 5648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5058
box 2028 5058 2228 5126
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4992
box 1832 4992 1900 5192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4830
box 2028 4830 2228 4898
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4764
box 1832 4764 1900 4964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5970
box 2028 5970 2228 6038
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5904
box 1832 5904 1900 6104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5286
box 2028 5286 2228 5354
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5220
box 1832 5220 1900 5420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5742
box 2028 5742 2228 5810
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5676
box 1832 5676 1900 5876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5514
box 2028 5514 2228 5582
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5448
box 1832 5448 1900 5648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5058
box 2028 5058 2228 5126
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4992
box 1832 4992 1900 5192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4830
box 2028 4830 2228 4898
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4764
box 1832 4764 1900 4964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5970
box 2028 5970 2228 6038
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5904
box 1832 5904 1900 6104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5286
box 2028 5286 2228 5354
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5220
box 1832 5220 1900 5420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5742
box 2028 5742 2228 5810
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5676
box 1832 5676 1900 5876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5514
box 2028 5514 2228 5582
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5448
box 1832 5448 1900 5648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5058
box 2028 5058 2228 5126
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4992
box 1832 4992 1900 5192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4830
box 2028 4830 2228 4898
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4764
box 1832 4764 1900 4964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5970
box 2028 5970 2228 6038
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5904
box 1832 5904 1900 6104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5286
box 2028 5286 2228 5354
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5220
box 1832 5220 1900 5420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5742
box 2028 5742 2228 5810
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5676
box 1832 5676 1900 5876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5514
box 2028 5514 2228 5582
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5448
box 1832 5448 1900 5648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5058
box 2028 5058 2228 5126
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4992
box 1832 4992 1900 5192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11006
box 2028 11006 2228 11074
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10940
box 1832 10940 1900 11140
use cut_M1M3_2x1 
transform 1 0 2028 0 1 12146
box 2028 12146 2228 12214
use cut_M2M3_1x2 
transform 1 0 1832 0 1 12080
box 1832 12080 1900 12280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11462
box 2028 11462 2228 11530
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11396
box 1832 11396 1900 11596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11918
box 2028 11918 2228 11986
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11852
box 1832 11852 1900 12052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11690
box 2028 11690 2228 11758
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11624
box 1832 11624 1900 11824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11234
box 2028 11234 2228 11302
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11168
box 1832 11168 1900 11368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11006
box 2028 11006 2228 11074
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10940
box 1832 10940 1900 11140
use cut_M1M3_2x1 
transform 1 0 2028 0 1 12146
box 2028 12146 2228 12214
use cut_M2M3_1x2 
transform 1 0 1832 0 1 12080
box 1832 12080 1900 12280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11462
box 2028 11462 2228 11530
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11396
box 1832 11396 1900 11596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11918
box 2028 11918 2228 11986
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11852
box 1832 11852 1900 12052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11690
box 2028 11690 2228 11758
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11624
box 1832 11624 1900 11824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11234
box 2028 11234 2228 11302
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11168
box 1832 11168 1900 11368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11006
box 2028 11006 2228 11074
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10940
box 1832 10940 1900 11140
use cut_M1M3_2x1 
transform 1 0 2028 0 1 12146
box 2028 12146 2228 12214
use cut_M2M3_1x2 
transform 1 0 1832 0 1 12080
box 1832 12080 1900 12280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11462
box 2028 11462 2228 11530
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11396
box 1832 11396 1900 11596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11918
box 2028 11918 2228 11986
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11852
box 1832 11852 1900 12052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11690
box 2028 11690 2228 11758
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11624
box 1832 11624 1900 11824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11234
box 2028 11234 2228 11302
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11168
box 1832 11168 1900 11368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11006
box 2028 11006 2228 11074
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10940
box 1832 10940 1900 11140
use cut_M1M3_2x1 
transform 1 0 2028 0 1 12146
box 2028 12146 2228 12214
use cut_M2M3_1x2 
transform 1 0 1832 0 1 12080
box 1832 12080 1900 12280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11462
box 2028 11462 2228 11530
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11396
box 1832 11396 1900 11596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11918
box 2028 11918 2228 11986
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11852
box 1832 11852 1900 12052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11690
box 2028 11690 2228 11758
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11624
box 1832 11624 1900 11824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11234
box 2028 11234 2228 11302
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11168
box 1832 11168 1900 11368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11006
box 2028 11006 2228 11074
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10940
box 1832 10940 1900 11140
use cut_M1M3_2x1 
transform 1 0 2028 0 1 12146
box 2028 12146 2228 12214
use cut_M2M3_1x2 
transform 1 0 1832 0 1 12080
box 1832 12080 1900 12280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11462
box 2028 11462 2228 11530
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11396
box 1832 11396 1900 11596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11918
box 2028 11918 2228 11986
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11852
box 1832 11852 1900 12052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11690
box 2028 11690 2228 11758
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11624
box 1832 11624 1900 11824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11234
box 2028 11234 2228 11302
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11168
box 1832 11168 1900 11368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11006
box 2028 11006 2228 11074
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10940
box 1832 10940 1900 11140
use cut_M1M3_2x1 
transform 1 0 2028 0 1 12146
box 2028 12146 2228 12214
use cut_M2M3_1x2 
transform 1 0 1832 0 1 12080
box 1832 12080 1900 12280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11462
box 2028 11462 2228 11530
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11396
box 1832 11396 1900 11596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11918
box 2028 11918 2228 11986
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11852
box 1832 11852 1900 12052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11690
box 2028 11690 2228 11758
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11624
box 1832 11624 1900 11824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11234
box 2028 11234 2228 11302
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11168
box 1832 11168 1900 11368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 198
box 2028 198 2228 266
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1338
box 2028 1338 2228 1406
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1272
box 1676 1272 1744 1472
use cut_M1M3_2x1 
transform 1 0 2028 0 1 654
box 2028 654 2228 722
use cut_M2M3_1x2 
transform 1 0 1676 0 1 588
box 1676 588 1744 788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1110
box 2028 1110 2228 1178
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1044
box 1676 1044 1744 1244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 882
box 2028 882 2228 950
use cut_M2M3_1x2 
transform 1 0 1676 0 1 816
box 1676 816 1744 1016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 426
box 2028 426 2228 494
use cut_M2M3_1x2 
transform 1 0 1676 0 1 360
box 1676 360 1744 560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 198
box 2028 198 2228 266
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1338
box 2028 1338 2228 1406
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1272
box 1676 1272 1744 1472
use cut_M1M3_2x1 
transform 1 0 2028 0 1 654
box 2028 654 2228 722
use cut_M2M3_1x2 
transform 1 0 1676 0 1 588
box 1676 588 1744 788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1110
box 2028 1110 2228 1178
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1044
box 1676 1044 1744 1244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 882
box 2028 882 2228 950
use cut_M2M3_1x2 
transform 1 0 1676 0 1 816
box 1676 816 1744 1016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 426
box 2028 426 2228 494
use cut_M2M3_1x2 
transform 1 0 1676 0 1 360
box 1676 360 1744 560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 198
box 2028 198 2228 266
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1338
box 2028 1338 2228 1406
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1272
box 1676 1272 1744 1472
use cut_M1M3_2x1 
transform 1 0 2028 0 1 654
box 2028 654 2228 722
use cut_M2M3_1x2 
transform 1 0 1676 0 1 588
box 1676 588 1744 788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1110
box 2028 1110 2228 1178
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1044
box 1676 1044 1744 1244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 882
box 2028 882 2228 950
use cut_M2M3_1x2 
transform 1 0 1676 0 1 816
box 1676 816 1744 1016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 426
box 2028 426 2228 494
use cut_M2M3_1x2 
transform 1 0 1676 0 1 360
box 1676 360 1744 560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 198
box 2028 198 2228 266
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1338
box 2028 1338 2228 1406
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1272
box 1676 1272 1744 1472
use cut_M1M3_2x1 
transform 1 0 2028 0 1 654
box 2028 654 2228 722
use cut_M2M3_1x2 
transform 1 0 1676 0 1 588
box 1676 588 1744 788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1110
box 2028 1110 2228 1178
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1044
box 1676 1044 1744 1244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 882
box 2028 882 2228 950
use cut_M2M3_1x2 
transform 1 0 1676 0 1 816
box 1676 816 1744 1016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 426
box 2028 426 2228 494
use cut_M2M3_1x2 
transform 1 0 1676 0 1 360
box 1676 360 1744 560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 198
box 2028 198 2228 266
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1338
box 2028 1338 2228 1406
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1272
box 1676 1272 1744 1472
use cut_M1M3_2x1 
transform 1 0 2028 0 1 654
box 2028 654 2228 722
use cut_M2M3_1x2 
transform 1 0 1676 0 1 588
box 1676 588 1744 788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1110
box 2028 1110 2228 1178
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1044
box 1676 1044 1744 1244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 882
box 2028 882 2228 950
use cut_M2M3_1x2 
transform 1 0 1676 0 1 816
box 1676 816 1744 1016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 426
box 2028 426 2228 494
use cut_M2M3_1x2 
transform 1 0 1676 0 1 360
box 1676 360 1744 560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 198
box 2028 198 2228 266
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1338
box 2028 1338 2228 1406
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1272
box 1676 1272 1744 1472
use cut_M1M3_2x1 
transform 1 0 2028 0 1 654
box 2028 654 2228 722
use cut_M2M3_1x2 
transform 1 0 1676 0 1 588
box 1676 588 1744 788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1110
box 2028 1110 2228 1178
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1044
box 1676 1044 1744 1244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 882
box 2028 882 2228 950
use cut_M2M3_1x2 
transform 1 0 1676 0 1 816
box 1676 816 1744 1016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 426
box 2028 426 2228 494
use cut_M2M3_1x2 
transform 1 0 1676 0 1 360
box 1676 360 1744 560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6374
box 2028 6374 2228 6442
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6308
box 1676 6308 1744 6508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7514
box 2028 7514 2228 7582
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7448
box 1676 7448 1744 7648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6830
box 2028 6830 2228 6898
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6764
box 1676 6764 1744 6964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7286
box 2028 7286 2228 7354
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7220
box 1676 7220 1744 7420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7058
box 2028 7058 2228 7126
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6992
box 1676 6992 1744 7192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6602
box 2028 6602 2228 6670
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6536
box 1676 6536 1744 6736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6374
box 2028 6374 2228 6442
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6308
box 1676 6308 1744 6508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7514
box 2028 7514 2228 7582
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7448
box 1676 7448 1744 7648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6830
box 2028 6830 2228 6898
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6764
box 1676 6764 1744 6964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7286
box 2028 7286 2228 7354
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7220
box 1676 7220 1744 7420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7058
box 2028 7058 2228 7126
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6992
box 1676 6992 1744 7192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6602
box 2028 6602 2228 6670
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6536
box 1676 6536 1744 6736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6374
box 2028 6374 2228 6442
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6308
box 1676 6308 1744 6508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7514
box 2028 7514 2228 7582
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7448
box 1676 7448 1744 7648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6830
box 2028 6830 2228 6898
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6764
box 1676 6764 1744 6964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7286
box 2028 7286 2228 7354
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7220
box 1676 7220 1744 7420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7058
box 2028 7058 2228 7126
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6992
box 1676 6992 1744 7192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6602
box 2028 6602 2228 6670
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6536
box 1676 6536 1744 6736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6374
box 2028 6374 2228 6442
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6308
box 1676 6308 1744 6508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7514
box 2028 7514 2228 7582
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7448
box 1676 7448 1744 7648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6830
box 2028 6830 2228 6898
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6764
box 1676 6764 1744 6964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7286
box 2028 7286 2228 7354
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7220
box 1676 7220 1744 7420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7058
box 2028 7058 2228 7126
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6992
box 1676 6992 1744 7192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6602
box 2028 6602 2228 6670
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6536
box 1676 6536 1744 6736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6374
box 2028 6374 2228 6442
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6308
box 1676 6308 1744 6508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7514
box 2028 7514 2228 7582
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7448
box 1676 7448 1744 7648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6830
box 2028 6830 2228 6898
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6764
box 1676 6764 1744 6964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7286
box 2028 7286 2228 7354
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7220
box 1676 7220 1744 7420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7058
box 2028 7058 2228 7126
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6992
box 1676 6992 1744 7192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6602
box 2028 6602 2228 6670
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6536
box 1676 6536 1744 6736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6374
box 2028 6374 2228 6442
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6308
box 1676 6308 1744 6508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7514
box 2028 7514 2228 7582
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7448
box 1676 7448 1744 7648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6830
box 2028 6830 2228 6898
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6764
box 1676 6764 1744 6964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7286
box 2028 7286 2228 7354
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7220
box 1676 7220 1744 7420
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7058
box 2028 7058 2228 7126
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6992
box 1676 6992 1744 7192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6602
box 2028 6602 2228 6670
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6536
box 1676 6536 1744 6736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9462
box 2028 9462 2228 9530
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9396
box 1520 9396 1588 9596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10602
box 2028 10602 2228 10670
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10536
box 1520 10536 1588 10736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9918
box 2028 9918 2228 9986
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9852
box 1520 9852 1588 10052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10374
box 2028 10374 2228 10442
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10308
box 1520 10308 1588 10508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10146
box 2028 10146 2228 10214
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10080
box 1520 10080 1588 10280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9690
box 2028 9690 2228 9758
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9624
box 1520 9624 1588 9824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9462
box 2028 9462 2228 9530
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9396
box 1520 9396 1588 9596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10602
box 2028 10602 2228 10670
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10536
box 1520 10536 1588 10736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9918
box 2028 9918 2228 9986
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9852
box 1520 9852 1588 10052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10374
box 2028 10374 2228 10442
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10308
box 1520 10308 1588 10508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10146
box 2028 10146 2228 10214
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10080
box 1520 10080 1588 10280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9690
box 2028 9690 2228 9758
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9624
box 1520 9624 1588 9824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9462
box 2028 9462 2228 9530
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9396
box 1520 9396 1588 9596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10602
box 2028 10602 2228 10670
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10536
box 1520 10536 1588 10736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9918
box 2028 9918 2228 9986
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9852
box 1520 9852 1588 10052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10374
box 2028 10374 2228 10442
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10308
box 1520 10308 1588 10508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10146
box 2028 10146 2228 10214
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10080
box 1520 10080 1588 10280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9690
box 2028 9690 2228 9758
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9624
box 1520 9624 1588 9824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9462
box 2028 9462 2228 9530
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9396
box 1520 9396 1588 9596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10602
box 2028 10602 2228 10670
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10536
box 1520 10536 1588 10736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9918
box 2028 9918 2228 9986
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9852
box 1520 9852 1588 10052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10374
box 2028 10374 2228 10442
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10308
box 1520 10308 1588 10508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10146
box 2028 10146 2228 10214
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10080
box 1520 10080 1588 10280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9690
box 2028 9690 2228 9758
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9624
box 1520 9624 1588 9824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9462
box 2028 9462 2228 9530
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9396
box 1520 9396 1588 9596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10602
box 2028 10602 2228 10670
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10536
box 1520 10536 1588 10736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9918
box 2028 9918 2228 9986
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9852
box 1520 9852 1588 10052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10374
box 2028 10374 2228 10442
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10308
box 1520 10308 1588 10508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10146
box 2028 10146 2228 10214
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10080
box 1520 10080 1588 10280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9690
box 2028 9690 2228 9758
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9624
box 1520 9624 1588 9824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9462
box 2028 9462 2228 9530
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9396
box 1520 9396 1588 9596
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10602
box 2028 10602 2228 10670
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10536
box 1520 10536 1588 10736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9918
box 2028 9918 2228 9986
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9852
box 1520 9852 1588 10052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10374
box 2028 10374 2228 10442
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10308
box 1520 10308 1588 10508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10146
box 2028 10146 2228 10214
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10080
box 1520 10080 1588 10280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9690
box 2028 9690 2228 9758
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9624
box 1520 9624 1588 9824
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1742
box 2028 1742 2228 1810
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1676
box 1364 1676 1432 1876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2882
box 2028 2882 2228 2950
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2816
box 1364 2816 1432 3016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2198
box 2028 2198 2228 2266
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2132
box 1364 2132 1432 2332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2654
box 2028 2654 2228 2722
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2588
box 1364 2588 1432 2788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2426
box 2028 2426 2228 2494
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2360
box 1364 2360 1432 2560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1970
box 2028 1970 2228 2038
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1904
box 1364 1904 1432 2104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1742
box 2028 1742 2228 1810
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1676
box 1364 1676 1432 1876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2882
box 2028 2882 2228 2950
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2816
box 1364 2816 1432 3016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2198
box 2028 2198 2228 2266
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2132
box 1364 2132 1432 2332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2654
box 2028 2654 2228 2722
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2588
box 1364 2588 1432 2788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2426
box 2028 2426 2228 2494
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2360
box 1364 2360 1432 2560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1970
box 2028 1970 2228 2038
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1904
box 1364 1904 1432 2104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1742
box 2028 1742 2228 1810
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1676
box 1364 1676 1432 1876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2882
box 2028 2882 2228 2950
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2816
box 1364 2816 1432 3016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2198
box 2028 2198 2228 2266
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2132
box 1364 2132 1432 2332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2654
box 2028 2654 2228 2722
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2588
box 1364 2588 1432 2788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2426
box 2028 2426 2228 2494
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2360
box 1364 2360 1432 2560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1970
box 2028 1970 2228 2038
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1904
box 1364 1904 1432 2104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1742
box 2028 1742 2228 1810
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1676
box 1364 1676 1432 1876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2882
box 2028 2882 2228 2950
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2816
box 1364 2816 1432 3016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2198
box 2028 2198 2228 2266
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2132
box 1364 2132 1432 2332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2654
box 2028 2654 2228 2722
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2588
box 1364 2588 1432 2788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2426
box 2028 2426 2228 2494
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2360
box 1364 2360 1432 2560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1970
box 2028 1970 2228 2038
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1904
box 1364 1904 1432 2104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1742
box 2028 1742 2228 1810
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1676
box 1364 1676 1432 1876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2882
box 2028 2882 2228 2950
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2816
box 1364 2816 1432 3016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2198
box 2028 2198 2228 2266
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2132
box 1364 2132 1432 2332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2654
box 2028 2654 2228 2722
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2588
box 1364 2588 1432 2788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2426
box 2028 2426 2228 2494
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2360
box 1364 2360 1432 2560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1970
box 2028 1970 2228 2038
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1904
box 1364 1904 1432 2104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1742
box 2028 1742 2228 1810
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1676
box 1364 1676 1432 1876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2882
box 2028 2882 2228 2950
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2816
box 1364 2816 1432 3016
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2198
box 2028 2198 2228 2266
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2132
box 1364 2132 1432 2332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2654
box 2028 2654 2228 2722
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2588
box 1364 2588 1432 2788
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2426
box 2028 2426 2228 2494
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2360
box 1364 2360 1432 2560
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1970
box 2028 1970 2228 2038
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1904
box 1364 1904 1432 2104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 3514
box 2028 3514 2228 3582
use cut_M2M3_1x2 
transform 1 0 1208 0 1 3448
box 1208 3448 1276 3648
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8146
box 2028 8146 2228 8214
use cut_M2M3_1x2 
transform 1 0 1052 0 1 8080
box 1052 8080 1120 8280
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7918
box 2028 7918 2228 7986
use cut_M2M3_1x2 
transform 1 0 896 0 1 7852
box 896 7852 964 8052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9058
box 2028 9058 2228 9126
use cut_M2M3_1x2 
transform 1 0 896 0 1 8992
box 896 8992 964 9192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8374
box 2028 8374 2228 8442
use cut_M2M3_1x2 
transform 1 0 896 0 1 8308
box 896 8308 964 8508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8830
box 2028 8830 2228 8898
use cut_M2M3_1x2 
transform 1 0 896 0 1 8764
box 896 8764 964 8964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7918
box 2028 7918 2228 7986
use cut_M2M3_1x2 
transform 1 0 896 0 1 7852
box 896 7852 964 8052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9058
box 2028 9058 2228 9126
use cut_M2M3_1x2 
transform 1 0 896 0 1 8992
box 896 8992 964 9192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8374
box 2028 8374 2228 8442
use cut_M2M3_1x2 
transform 1 0 896 0 1 8308
box 896 8308 964 8508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8830
box 2028 8830 2228 8898
use cut_M2M3_1x2 
transform 1 0 896 0 1 8764
box 896 8764 964 8964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7918
box 2028 7918 2228 7986
use cut_M2M3_1x2 
transform 1 0 896 0 1 7852
box 896 7852 964 8052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9058
box 2028 9058 2228 9126
use cut_M2M3_1x2 
transform 1 0 896 0 1 8992
box 896 8992 964 9192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8374
box 2028 8374 2228 8442
use cut_M2M3_1x2 
transform 1 0 896 0 1 8308
box 896 8308 964 8508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8830
box 2028 8830 2228 8898
use cut_M2M3_1x2 
transform 1 0 896 0 1 8764
box 896 8764 964 8964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7918
box 2028 7918 2228 7986
use cut_M2M3_1x2 
transform 1 0 896 0 1 7852
box 896 7852 964 8052
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9058
box 2028 9058 2228 9126
use cut_M2M3_1x2 
transform 1 0 896 0 1 8992
box 896 8992 964 9192
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8374
box 2028 8374 2228 8442
use cut_M2M3_1x2 
transform 1 0 896 0 1 8308
box 896 8308 964 8508
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8830
box 2028 8830 2228 8898
use cut_M2M3_1x2 
transform 1 0 896 0 1 8764
box 896 8764 964 8964
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8602
box 2028 8602 2228 8670
use cut_M2M3_1x2 
transform 1 0 740 0 1 8536
box 740 8536 808 8736
use cut_M1M3_2x1 
transform 1 0 2028 0 1 3970
box 2028 3970 2228 4038
use cut_M2M3_1x2 
transform 1 0 584 0 1 3904
box 584 3904 652 4104
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4198
box 2028 4198 2228 4266
use cut_M2M3_1x2 
transform 1 0 428 0 1 4132
box 428 4132 496 4332
use cut_M1M3_2x1 
transform 1 0 2028 0 1 3742
box 2028 3742 2228 3810
use cut_M2M3_1x2 
transform 1 0 272 0 1 3676
box 272 3676 340 3876
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4426
box 2028 4426 2228 4494
use cut_M2M3_1x2 
transform 1 0 116 0 1 4360
box 116 4360 184 4560
use cut_M1M2_1x2 
transform 1 0 2356 0 1 3220
box 2356 3220 2424 3420
use cut_M1M2_1x2 
transform 1 0 2356 0 1 3220
box 2356 3220 2424 3420
<< labels >>
flabel m1 s 1836 4764 1896 12352 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew
flabel m1 s 1680 132 1740 12352 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew
flabel m1 s 1524 9396 1584 12352 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew
flabel m1 s 1368 1676 1428 12352 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew
flabel m1 s 1212 3448 1272 12352 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew
flabel m1 s 1056 8080 1116 12352 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew
flabel m1 s 900 7852 960 12352 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew
flabel m1 s 744 8536 804 12352 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew
flabel m1 s 588 3904 648 12352 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew
flabel m1 s 432 4132 492 12352 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew
flabel m1 s 276 3676 336 12352 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew
flabel m1 s 120 4360 180 12352 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew
flabel m1 s 2356 0 10936 68 0 FreeSans 400 0 0 0 AVSS
port 13 nsew
flabel m3 s 2356 10808 2424 12412 0 FreeSans 400 0 0 0 CTOP
port 14 nsew
<< end >>
