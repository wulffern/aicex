* NGSPICE file created from SUNTR_CAP_10.ext - technology: sky130A

.subckt SUNTR_CAP_10 A B
R0 A m3_2628_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R1 m3_252_308# B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
C0 A B 25.81fF
C1 B 0 5.39fF
C2 A 0 5.36fF
.ends
