magic
tech sky130A
magscale 1 2
timestamp 1660215182
<< checkpaint >>
rect -640 -640 3016 3500
<< locali >>
rect -640 -640 3016 -528
rect -640 -640 3016 -528
rect -640 -640 -528 3500
rect -640 3388 3016 3500
rect 2904 -640 3016 3500
rect -640 -640 3016 -528
rect 2106 2750 2430 2970
rect -54 2750 270 2970
<< ptapc >>
rect -612 -640 -532 -560
rect -532 -640 -452 -560
rect -452 -640 -372 -560
rect -372 -640 -292 -560
rect -292 -640 -212 -560
rect -212 -640 -132 -560
rect -132 -640 -52 -560
rect -52 -640 28 -560
rect 28 -640 108 -560
rect 108 -640 188 -560
rect 188 -640 268 -560
rect 268 -640 348 -560
rect 348 -640 428 -560
rect 428 -640 508 -560
rect 508 -640 588 -560
rect 588 -640 668 -560
rect 668 -640 748 -560
rect 748 -640 828 -560
rect 828 -640 908 -560
rect 908 -640 988 -560
rect 988 -640 1068 -560
rect 1068 -640 1148 -560
rect 1148 -640 1228 -560
rect 1228 -640 1308 -560
rect 1308 -640 1388 -560
rect 1388 -640 1468 -560
rect 1468 -640 1548 -560
rect 1548 -640 1628 -560
rect 1628 -640 1708 -560
rect 1708 -640 1788 -560
rect 1788 -640 1868 -560
rect 1868 -640 1948 -560
rect 1948 -640 2028 -560
rect 2028 -640 2108 -560
rect 2108 -640 2188 -560
rect 2188 -640 2268 -560
rect 2268 -640 2348 -560
rect 2348 -640 2428 -560
rect 2428 -640 2508 -560
rect 2508 -640 2588 -560
rect 2588 -640 2668 -560
rect 2668 -640 2748 -560
rect 2748 -640 2828 -560
rect 2828 -640 2908 -560
rect 2908 -640 2988 -560
rect -640 -610 -560 -530
rect -640 -530 -560 -450
rect -640 -450 -560 -370
rect -640 -370 -560 -290
rect -640 -290 -560 -210
rect -640 -210 -560 -130
rect -640 -130 -560 -50
rect -640 -50 -560 30
rect -640 30 -560 110
rect -640 110 -560 190
rect -640 190 -560 270
rect -640 270 -560 350
rect -640 350 -560 430
rect -640 430 -560 510
rect -640 510 -560 590
rect -640 590 -560 670
rect -640 670 -560 750
rect -640 750 -560 830
rect -640 830 -560 910
rect -640 910 -560 990
rect -640 990 -560 1070
rect -640 1070 -560 1150
rect -640 1150 -560 1230
rect -640 1230 -560 1310
rect -640 1310 -560 1390
rect -640 1390 -560 1470
rect -640 1470 -560 1550
rect -640 1550 -560 1630
rect -640 1630 -560 1710
rect -640 1710 -560 1790
rect -640 1790 -560 1870
rect -640 1870 -560 1950
rect -640 1950 -560 2030
rect -640 2030 -560 2110
rect -640 2110 -560 2190
rect -640 2190 -560 2270
rect -640 2270 -560 2350
rect -640 2350 -560 2430
rect -640 2430 -560 2510
rect -640 2510 -560 2590
rect -640 2590 -560 2670
rect -640 2670 -560 2750
rect -640 2750 -560 2830
rect -640 2830 -560 2910
rect -640 2910 -560 2990
rect -640 2990 -560 3070
rect -640 3070 -560 3150
rect -640 3150 -560 3230
rect -640 3230 -560 3310
rect -640 3310 -560 3390
rect -640 3390 -560 3470
rect -612 3388 -532 3468
rect -532 3388 -452 3468
rect -452 3388 -372 3468
rect -372 3388 -292 3468
rect -292 3388 -212 3468
rect -212 3388 -132 3468
rect -132 3388 -52 3468
rect -52 3388 28 3468
rect 28 3388 108 3468
rect 108 3388 188 3468
rect 188 3388 268 3468
rect 268 3388 348 3468
rect 348 3388 428 3468
rect 428 3388 508 3468
rect 508 3388 588 3468
rect 588 3388 668 3468
rect 668 3388 748 3468
rect 748 3388 828 3468
rect 828 3388 908 3468
rect 908 3388 988 3468
rect 988 3388 1068 3468
rect 1068 3388 1148 3468
rect 1148 3388 1228 3468
rect 1228 3388 1308 3468
rect 1308 3388 1388 3468
rect 1388 3388 1468 3468
rect 1468 3388 1548 3468
rect 1548 3388 1628 3468
rect 1628 3388 1708 3468
rect 1708 3388 1788 3468
rect 1788 3388 1868 3468
rect 1868 3388 1948 3468
rect 1948 3388 2028 3468
rect 2028 3388 2108 3468
rect 2108 3388 2188 3468
rect 2188 3388 2268 3468
rect 2268 3388 2348 3468
rect 2348 3388 2428 3468
rect 2428 3388 2508 3468
rect 2508 3388 2588 3468
rect 2588 3388 2668 3468
rect 2668 3388 2748 3468
rect 2748 3388 2828 3468
rect 2828 3388 2908 3468
rect 2908 3388 2988 3468
rect 2904 -610 2984 -530
rect 2904 -530 2984 -450
rect 2904 -450 2984 -370
rect 2904 -370 2984 -290
rect 2904 -290 2984 -210
rect 2904 -210 2984 -130
rect 2904 -130 2984 -50
rect 2904 -50 2984 30
rect 2904 30 2984 110
rect 2904 110 2984 190
rect 2904 190 2984 270
rect 2904 270 2984 350
rect 2904 350 2984 430
rect 2904 430 2984 510
rect 2904 510 2984 590
rect 2904 590 2984 670
rect 2904 670 2984 750
rect 2904 750 2984 830
rect 2904 830 2984 910
rect 2904 910 2984 990
rect 2904 990 2984 1070
rect 2904 1070 2984 1150
rect 2904 1150 2984 1230
rect 2904 1230 2984 1310
rect 2904 1310 2984 1390
rect 2904 1390 2984 1470
rect 2904 1470 2984 1550
rect 2904 1550 2984 1630
rect 2904 1630 2984 1710
rect 2904 1710 2984 1790
rect 2904 1790 2984 1870
rect 2904 1870 2984 1950
rect 2904 1950 2984 2030
rect 2904 2030 2984 2110
rect 2904 2110 2984 2190
rect 2904 2190 2984 2270
rect 2904 2270 2984 2350
rect 2904 2350 2984 2430
rect 2904 2430 2984 2510
rect 2904 2510 2984 2590
rect 2904 2590 2984 2670
rect 2904 2670 2984 2750
rect 2904 2750 2984 2830
rect 2904 2830 2984 2910
rect 2904 2910 2984 2990
rect 2904 2990 2984 3070
rect 2904 3070 2984 3150
rect 2904 3150 2984 3230
rect 2904 3230 2984 3310
rect 2904 3310 2984 3390
rect 2904 3390 2984 3470
<< ptap >>
rect -640 -640 3016 -528
rect -640 -640 -528 3500
rect -640 3388 3016 3500
rect 2904 -640 3016 3500
use SUNTR_RES100 XA1
transform 1 0 0 0 1 0
box 0 0 2376 2860
<< labels >>
flabel locali s -640 -640 3016 -528 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 2106 2750 2430 2970 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s -54 2750 270 2970 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
