magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 2240
<< locali >>
rect 690 210 750 2030
rect 720 210 874 270
rect 874 50 1380 110
rect 874 50 934 270
rect 330 450 390 1790
rect 1710 450 1770 2110
rect 1350 210 1410 2190
rect 630 2130 1470 2190
rect 1380 2130 1534 2190
rect 1534 2050 1740 2110
rect 1534 2050 1594 2190
rect 690 210 750 430
rect 690 530 750 750
rect 690 850 750 1070
rect 690 1170 750 1390
rect 690 1490 750 1710
rect 690 1810 750 2030
rect 1350 210 1410 430
rect 1350 530 1410 750
rect 1350 850 1410 1070
rect 1350 1170 1410 1390
rect 1350 1490 1410 1710
rect 1350 1810 1410 2030
rect 2010 120 2190 200
rect -90 120 90 200
rect 270 2050 450 2110
rect 270 130 450 190
rect 270 450 450 510
<< poly >>
rect 270 142 1830 178
<< m3 >>
rect 1290 0 1474 2240
rect 630 0 814 2240
rect 1290 0 1474 2240
rect 630 0 814 2240
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1050 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1050 1280
use NCHDL MN4
transform 1 0 0 0 1 1280
box 0 1280 1050 1600
use NCHDL MN5
transform 1 0 0 0 1 1600
box 0 1600 1050 1920
use NCHDL MN6
transform 1 0 0 0 1 1920
box 0 1920 1050 2240
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1_DMY
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL MP2_DMY
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use PCHDL MP3_DMY
transform 1 0 1050 0 1 960
box 1050 960 2100 1280
use PCHDL MP4_DMY
transform 1 0 1050 0 1 1280
box 1050 1280 2100 1600
use PCHDL MP5_DMY
transform 1 0 1050 0 1 1600
box 1050 1600 2100 1920
use PCHDL MP6_DMY
transform 1 0 1050 0 1 1920
box 1050 1920 2100 2240
use cut_M1M4_2x1 
transform 1 0 1290 0 1 210
box 1290 210 1474 278
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
<< labels >>
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 270 2050 450 2110 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 CKN
port 4 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 CI
port 5 nsew
flabel m3 s 1290 0 1474 2240 0 FreeSans 400 0 0 0 AVDD
port 6 nsew
flabel m3 s 630 0 814 2240 0 FreeSans 400 0 0 0 AVSS
port 7 nsew
<< end >>
