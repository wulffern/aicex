magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect -2028 -1560 24252 38534
<< m3 >>
rect 8580 17384 22702 17444
rect 8580 17724 22702 17784
rect 20562 18056 20622 24704
rect 20790 18056 20850 31744
rect 4722 18124 4782 27900
rect 5438 18294 5498 27900
rect 8682 18464 8742 27900
rect 1478 18634 1538 27900
rect 12078 18804 12138 27922
rect 16038 18974 16098 27922
rect 10078 19144 10138 27922
rect 14038 19314 14098 27922
rect 2158 19484 2218 27922
rect 6118 19654 6178 27922
rect 4158 19824 4218 27922
rect 8118 19994 8178 27922
rect 2294 20164 2354 29202
rect 7982 20334 8042 29202
rect 6254 20504 6314 29202
rect 4022 20674 4082 29202
rect 10350 20844 10410 30482
rect 11806 21014 11866 30482
rect 14310 21184 14370 30482
rect 7846 21354 7906 30482
rect 3886 21524 3946 30482
rect 2430 21694 2490 30482
rect 15766 21864 15826 30482
rect 6390 22034 6450 30482
rect 1842 22654 2026 37334
rect 4358 22654 4542 37334
rect 5802 22654 5986 37334
rect 8318 22654 8502 37334
rect 9762 22654 9946 37334
rect 12278 22654 12462 37334
rect 13722 22654 13906 37334
rect 16238 22654 16422 37334
rect 17682 22654 17866 37334
rect 20198 22654 20382 37334
rect 9158 -600 9342 4800
rect 12882 -600 13066 4800
rect 2382 22654 2566 37934
rect 3818 22654 4002 37934
rect 6342 22654 6526 37934
rect 7778 22654 7962 37934
rect 10302 22654 10486 37934
rect 11738 22654 11922 37934
rect 14262 22654 14446 37934
rect 15698 22654 15882 37934
rect 18222 22654 18406 37934
rect 19658 22654 19842 37934
rect 8618 -1200 8802 4800
rect 13422 -1200 13606 4800
rect 2862 27024 3046 38534
rect 3338 27024 3522 38534
rect 6822 27024 7006 38534
rect 7298 27024 7482 38534
rect 10782 27024 10966 38534
rect 11258 27024 11442 38534
rect 14742 27024 14926 38534
rect 15218 27024 15402 38534
rect 18702 27024 18886 38534
rect 9776 -1560 9836 3154
rect 12388 -1560 12448 3154
rect 10194 1170 10392 1230
rect 8614 4970 10194 5030
rect 11832 1170 11970 1230
rect 11970 4970 13606 5030
rect 10392 1170 10530 1230
rect 10530 2450 11832 2510
rect 10530 1170 10590 2518
<< m2 >>
rect 13572 16934 13632 17452
rect 8580 16934 8640 17792
rect 4722 18064 12816 18124
rect 5438 18234 12504 18294
rect 8682 18404 12192 18464
rect 1478 18574 13128 18634
rect 10496 18744 12138 18804
rect 10808 18914 16098 18974
rect 10078 19084 10400 19144
rect 10652 19254 14098 19314
rect 2158 19424 9152 19484
rect 6118 19594 9776 19654
rect 4158 19764 9464 19824
rect 8118 19934 10088 19994
rect 2294 20104 9308 20164
rect 7982 20274 10244 20334
rect 6254 20444 9932 20504
rect 4022 20614 9620 20674
rect 10350 20784 11880 20844
rect 11664 20954 11866 21014
rect 11508 21124 14370 21184
rect 7846 21294 12036 21354
rect 3886 21464 12660 21524
rect 2430 21634 12972 21694
rect 11352 21804 15826 21864
rect 6390 21974 12348 22034
rect 2382 35374 2658 35434
rect 2658 34836 4722 34896
rect 4662 34836 4722 35004
rect 2658 34836 2718 35446
rect 6342 35374 6618 35434
rect 6618 34836 8682 34896
rect 8622 34836 8682 35004
rect 6618 34836 6678 35446
rect 10302 35374 10578 35434
rect 10578 34836 12642 34896
rect 12582 34836 12642 35004
rect 10578 34836 10638 35446
rect 14262 35374 14538 35434
rect 14538 34836 16602 34896
rect 16542 34836 16602 35004
rect 14538 34836 14598 35446
rect 1482 31956 17502 32016
rect 1422 31956 1482 32124
rect 4662 31956 4722 32124
rect 5382 31956 5442 32124
rect 8622 31956 8682 32124
rect 9342 31956 9402 32124
rect 12582 31956 12642 32124
rect 13302 31956 13362 32124
rect 16542 31956 16602 32124
rect 17262 31956 17322 32124
rect 2378 23340 2658 23400
rect 2658 22992 4722 23052
rect 4662 22992 4722 23168
rect 2658 22992 2718 23400
rect 6338 23340 6618 23400
rect 6618 22992 8682 23052
rect 8622 22992 8682 23168
rect 6618 22992 6678 23400
rect 10298 23340 10578 23400
rect 10578 22992 12642 23052
rect 12582 22992 12642 23168
rect 10578 22992 10638 23400
rect 14258 23340 14538 23400
rect 14538 22992 16602 23052
rect 16542 22992 16602 23168
rect 14538 22992 14598 23400
rect 18218 23340 18498 23400
rect 18498 23340 18558 23400
rect 3822 23340 4102 23400
rect 4102 23340 4162 23448
rect 4102 23448 5438 23508
rect 5378 23100 5438 23508
rect 7782 23340 8062 23400
rect 8062 23340 8122 23448
rect 8062 23448 9398 23508
rect 9338 23100 9398 23508
rect 11742 23340 12022 23400
rect 12022 23340 12082 23448
rect 12022 23448 13358 23508
rect 13298 23100 13358 23508
rect 15702 23340 15982 23400
rect 15982 23340 16042 23448
rect 15982 23448 17318 23508
rect 17258 23100 17318 23508
rect 1478 25024 17502 25084
rect 1418 24700 1478 25084
rect 4662 24700 4722 25084
rect 5378 24700 5438 25084
rect 8622 24700 8682 25084
rect 9338 24700 9398 25084
rect 12582 24700 12642 25084
rect 13298 24700 13358 25084
rect 16542 24700 16602 25084
rect 17258 24700 17318 25084
rect 1482 25348 17502 25408
rect 1422 25348 1482 25724
rect 4662 25348 4722 25724
rect 5382 25348 5442 25724
rect 8622 25348 8682 25724
rect 9342 25348 9402 25724
rect 12582 25348 12642 25724
rect 13302 25348 13362 25724
rect 16542 25348 16602 25724
rect 17262 25348 17322 25724
rect 2742 26304 1662 26364
rect 2742 26304 2922 26364
rect 2742 26304 3642 26364
rect 2742 26304 6882 26364
rect 2742 26304 7602 26364
rect 2742 26304 10842 26364
rect 2742 26304 11562 26364
rect 2742 26304 14802 26364
rect 2742 26304 15522 26364
rect 2742 26304 18762 26364
rect 20094 27694 20292 27754
rect 17442 24760 20094 24820
rect 20094 24760 20154 27766
rect 17410 24700 17502 24760
rect 19554 28974 19752 29034
rect 17442 25724 19554 25784
rect 19554 25724 19614 29046
rect 17412 25664 17502 25724
rect 19392 35584 19530 35644
rect 17412 32704 19530 32764
rect 19530 32704 19590 35652
rect 19194 36224 19392 36284
rect 18312 35374 19194 35434
rect 19194 35374 19254 36292
rect 10392 2450 10530 2510
rect 10530 1170 11832 1230
rect 10530 1170 10590 2518
rect 1482 26304 2922 26364
<< m4 >>
rect 20562 17724 20622 18056
rect 20790 17384 20850 18056
rect 10194 1170 10254 5030
rect 11970 1170 12030 5030
<< m1 >>
rect 12756 16874 12816 18064
rect 12444 16874 12504 18234
rect 12132 16874 12192 18404
rect 13068 16874 13128 18574
rect 10496 16874 10556 18744
rect 10808 16874 10868 18914
rect 10340 16874 10400 19084
rect 10652 16874 10712 19254
rect 9092 16874 9152 19424
rect 9716 16874 9776 19594
rect 9404 16874 9464 19764
rect 10028 16874 10088 19934
rect 9248 16874 9308 20104
rect 10184 16874 10244 20274
rect 9872 16874 9932 20444
rect 9560 16874 9620 20614
rect 11820 16874 11880 20784
rect 11664 16874 11724 20954
rect 11508 16874 11568 21124
rect 11976 16874 12036 21294
rect 12600 16874 12660 21464
rect 12912 16874 12972 21634
rect 11352 16874 11412 21804
rect 12288 16874 12348 21974
rect 9582 -1380 9642 510
rect 12582 -1380 12642 510
rect 1482 34944 -1968 35004
rect 3822 35344 4098 35404
rect 4098 34836 5442 34896
rect 5382 34836 5442 35004
rect 4098 34836 4158 35412
rect 7782 35344 8058 35404
rect 8058 34836 9402 34896
rect 9342 34836 9402 35004
rect 8058 34836 8118 35412
rect 11742 35344 12018 35404
rect 12018 34836 13362 34896
rect 13302 34836 13362 35004
rect 12018 34836 12078 35412
rect 15702 35344 15978 35404
rect 15978 34836 17322 34896
rect 17262 34836 17322 35004
rect 15978 34836 16038 35412
rect 19194 35904 19392 35964
rect 17772 33424 19194 33484
rect 19194 33424 19254 35972
rect -1248 4970 68 5030
rect -1248 6458 68 6518
rect -1248 7946 68 8006
rect -1248 9434 68 9494
rect -1248 10922 68 10982
rect -1248 12410 68 12470
rect -1248 13898 68 13958
rect -1248 15386 68 15446
rect 22152 4970 23472 5030
rect 22152 6458 23472 6518
rect 22152 7946 23472 8006
rect 22152 9434 23472 9494
rect 22152 10922 23472 10982
rect 22152 12410 23472 12470
rect 22152 13898 23472 13958
rect 22152 15386 23472 15446
<< locali >>
rect -1248 -600 23472 -416
rect -1248 37150 23472 37334
rect -1248 -600 -1064 37334
rect 23288 -600 23472 37334
rect -1848 -1200 24072 -1016
rect -1848 37750 24072 37934
rect -1848 -1200 -1664 37934
rect 23888 -1200 24072 37934
rect -1848 38350 24072 38534
rect -1848 -1380 24252 -1320
rect 24192 -1380 24252 38534
rect -2028 -1560 24252 -1500
rect -2028 -1560 -1968 38534
use SARBSSW_CV XB1
transform -1 0 11112 0 1 0
box 11112 0 22872 4800
use SARBSSW_CV XB2
transform 1 0 11112 0 1 0
box 11112 0 22872 4800
use CDAC8_CV XDAC1
transform -1 0 10988 0 1 4970
box 10988 4970 21860 16934
use CDAC8_CV XDAC2
transform 1 0 11232 0 1 4970
box 11232 4970 22104 16934
use SARDIGEX4_CV XA0
transform 1 0 1212 0 1 22654
box 1212 22654 3192 35774
use SARDIGEX4_CV XA1
transform -1 0 5172 0 1 22654
box 5172 22654 7152 35774
use SARDIGEX4_CV XA2
transform 1 0 5172 0 1 22654
box 5172 22654 7152 35774
use SARDIGEX4_CV XA3
transform -1 0 9132 0 1 22654
box 9132 22654 11112 35774
use SARDIGEX4_CV XA4
transform 1 0 9132 0 1 22654
box 9132 22654 11112 35774
use SARDIGEX4_CV XA5
transform -1 0 13092 0 1 22654
box 13092 22654 15072 35774
use SARDIGEX4_CV XA6
transform 1 0 13092 0 1 22654
box 13092 22654 15072 35774
use SARDIGEX4_CV XA7
transform -1 0 17052 0 1 22654
box 17052 22654 19032 35774
use SARDIGEX4_CV XA8
transform 1 0 17052 0 1 22654
box 17052 22654 19032 35774
use SARCMPX1_CV XA20
transform -1 0 21012 0 1 22654
box 21012 22654 22992 36734
use cut_M3M4_1x2 
transform 1 0 13572 0 1 16934
box 13572 16934 13640 17118
use cut_M3M4_2x1 
transform 1 0 13572 0 1 17384
box 13572 17384 13756 17452
use cut_M3M4_1x2 
transform 1 0 8580 0 1 16934
box 8580 16934 8648 17118
use cut_M3M4_2x1 
transform 1 0 8580 0 1 17724
box 8580 17724 8764 17792
use cut_M2M4_2x1 
transform 1 0 20562 0 1 24704
box 20562 24704 20746 24772
use cut_M4M5_2x1 
transform 1 0 20562 0 1 17724
box 20562 17724 20746 17792
use cut_M4M5_1x2 
transform 1 0 20562 0 1 18056
box 20562 18056 20630 18240
use cut_M3M4_2x1 
transform 1 0 20666 0 1 31744
box 20666 31744 20850 31812
use cut_M2M3_2x1 
transform 1 0 20562 0 1 31744
box 20562 31744 20746 31812
use cut_M4M5_2x1 
transform 1 0 20790 0 1 17384
box 20790 17384 20974 17452
use cut_M4M5_1x2 
transform 1 0 20790 0 1 18056
box 20790 18056 20858 18240
use cut_M3M4_1x2 
transform 1 0 4718 0 1 18002
box 4718 18002 4786 18186
use cut_M2M3_1x2 
transform 1 0 12752 0 1 18002
box 12752 18002 12820 18186
use cut_M3M4_1x2 
transform 1 0 5434 0 1 18172
box 5434 18172 5502 18356
use cut_M2M3_1x2 
transform 1 0 12440 0 1 18172
box 12440 18172 12508 18356
use cut_M3M4_1x2 
transform 1 0 8678 0 1 18342
box 8678 18342 8746 18526
use cut_M2M3_1x2 
transform 1 0 12128 0 1 18342
box 12128 18342 12196 18526
use cut_M3M4_1x2 
transform 1 0 1474 0 1 18512
box 1474 18512 1542 18696
use cut_M2M3_1x2 
transform 1 0 13064 0 1 18512
box 13064 18512 13132 18696
use cut_M3M4_1x2 
transform 1 0 12074 0 1 18682
box 12074 18682 12142 18866
use cut_M2M3_1x2 
transform 1 0 10492 0 1 18682
box 10492 18682 10560 18866
use cut_M3M4_1x2 
transform 1 0 16034 0 1 18852
box 16034 18852 16102 19036
use cut_M2M3_1x2 
transform 1 0 10804 0 1 18852
box 10804 18852 10872 19036
use cut_M3M4_1x2 
transform 1 0 10074 0 1 19022
box 10074 19022 10142 19206
use cut_M2M3_1x2 
transform 1 0 10336 0 1 19022
box 10336 19022 10404 19206
use cut_M3M4_1x2 
transform 1 0 14034 0 1 19192
box 14034 19192 14102 19376
use cut_M2M3_1x2 
transform 1 0 10648 0 1 19192
box 10648 19192 10716 19376
use cut_M3M4_1x2 
transform 1 0 2154 0 1 19362
box 2154 19362 2222 19546
use cut_M2M3_1x2 
transform 1 0 9088 0 1 19362
box 9088 19362 9156 19546
use cut_M3M4_1x2 
transform 1 0 6114 0 1 19532
box 6114 19532 6182 19716
use cut_M2M3_1x2 
transform 1 0 9712 0 1 19532
box 9712 19532 9780 19716
use cut_M3M4_1x2 
transform 1 0 4154 0 1 19702
box 4154 19702 4222 19886
use cut_M2M3_1x2 
transform 1 0 9400 0 1 19702
box 9400 19702 9468 19886
use cut_M3M4_1x2 
transform 1 0 8114 0 1 19872
box 8114 19872 8182 20056
use cut_M2M3_1x2 
transform 1 0 10024 0 1 19872
box 10024 19872 10092 20056
use cut_M3M4_1x2 
transform 1 0 2290 0 1 20042
box 2290 20042 2358 20226
use cut_M2M3_1x2 
transform 1 0 9244 0 1 20042
box 9244 20042 9312 20226
use cut_M3M4_1x2 
transform 1 0 7978 0 1 20212
box 7978 20212 8046 20396
use cut_M2M3_1x2 
transform 1 0 10180 0 1 20212
box 10180 20212 10248 20396
use cut_M3M4_1x2 
transform 1 0 6250 0 1 20382
box 6250 20382 6318 20566
use cut_M2M3_1x2 
transform 1 0 9868 0 1 20382
box 9868 20382 9936 20566
use cut_M3M4_1x2 
transform 1 0 4018 0 1 20552
box 4018 20552 4086 20736
use cut_M2M3_1x2 
transform 1 0 9556 0 1 20552
box 9556 20552 9624 20736
use cut_M3M4_1x2 
transform 1 0 10346 0 1 20722
box 10346 20722 10414 20906
use cut_M2M3_1x2 
transform 1 0 11816 0 1 20722
box 11816 20722 11884 20906
use cut_M3M4_1x2 
transform 1 0 11802 0 1 20892
box 11802 20892 11870 21076
use cut_M2M3_1x2 
transform 1 0 11660 0 1 20892
box 11660 20892 11728 21076
use cut_M3M4_1x2 
transform 1 0 14306 0 1 21062
box 14306 21062 14374 21246
use cut_M2M3_1x2 
transform 1 0 11504 0 1 21062
box 11504 21062 11572 21246
use cut_M3M4_1x2 
transform 1 0 7842 0 1 21232
box 7842 21232 7910 21416
use cut_M2M3_1x2 
transform 1 0 11972 0 1 21232
box 11972 21232 12040 21416
use cut_M3M4_1x2 
transform 1 0 3882 0 1 21402
box 3882 21402 3950 21586
use cut_M2M3_1x2 
transform 1 0 12596 0 1 21402
box 12596 21402 12664 21586
use cut_M3M4_1x2 
transform 1 0 2426 0 1 21572
box 2426 21572 2494 21756
use cut_M2M3_1x2 
transform 1 0 12908 0 1 21572
box 12908 21572 12976 21756
use cut_M3M4_1x2 
transform 1 0 15762 0 1 21742
box 15762 21742 15830 21926
use cut_M2M3_1x2 
transform 1 0 11348 0 1 21742
box 11348 21742 11416 21926
use cut_M3M4_1x2 
transform 1 0 6386 0 1 21912
box 6386 21912 6454 22096
use cut_M2M3_1x2 
transform 1 0 12284 0 1 21912
box 12284 21912 12352 22096
use cut_M1M4_2x2 
transform 1 0 1842 0 1 37150
box 1842 37150 2026 37334
use cut_M1M4_2x2 
transform 1 0 4358 0 1 37150
box 4358 37150 4542 37334
use cut_M1M4_2x2 
transform 1 0 5802 0 1 37150
box 5802 37150 5986 37334
use cut_M1M4_2x2 
transform 1 0 8318 0 1 37150
box 8318 37150 8502 37334
use cut_M1M4_2x2 
transform 1 0 9762 0 1 37150
box 9762 37150 9946 37334
use cut_M1M4_2x2 
transform 1 0 12278 0 1 37150
box 12278 37150 12462 37334
use cut_M1M4_2x2 
transform 1 0 13722 0 1 37150
box 13722 37150 13906 37334
use cut_M1M4_2x2 
transform 1 0 16238 0 1 37150
box 16238 37150 16422 37334
use cut_M1M4_2x2 
transform 1 0 17682 0 1 37150
box 17682 37150 17866 37334
use cut_M1M4_2x2 
transform 1 0 20198 0 1 37150
box 20198 37150 20382 37334
use cut_M1M4_2x2 
transform 1 0 9158 0 1 -600
box 9158 -600 9342 -416
use cut_M1M4_2x2 
transform 1 0 12882 0 1 -600
box 12882 -600 13066 -416
use cut_M1M4_2x2 
transform 1 0 2382 0 1 37750
box 2382 37750 2566 37934
use cut_M1M4_2x2 
transform 1 0 3818 0 1 37750
box 3818 37750 4002 37934
use cut_M1M4_2x2 
transform 1 0 6342 0 1 37750
box 6342 37750 6526 37934
use cut_M1M4_2x2 
transform 1 0 7778 0 1 37750
box 7778 37750 7962 37934
use cut_M1M4_2x2 
transform 1 0 10302 0 1 37750
box 10302 37750 10486 37934
use cut_M1M4_2x2 
transform 1 0 11738 0 1 37750
box 11738 37750 11922 37934
use cut_M1M4_2x2 
transform 1 0 14262 0 1 37750
box 14262 37750 14446 37934
use cut_M1M4_2x2 
transform 1 0 15698 0 1 37750
box 15698 37750 15882 37934
use cut_M1M4_2x2 
transform 1 0 18222 0 1 37750
box 18222 37750 18406 37934
use cut_M1M4_2x2 
transform 1 0 19658 0 1 37750
box 19658 37750 19842 37934
use cut_M1M4_2x2 
transform 1 0 8618 0 1 -1200
box 8618 -1200 8802 -1016
use cut_M1M4_2x2 
transform 1 0 13422 0 1 -1200
box 13422 -1200 13606 -1016
use cut_M1M4_2x2 
transform 1 0 2862 0 1 38350
box 2862 38350 3046 38534
use cut_M1M4_2x2 
transform 1 0 3338 0 1 38350
box 3338 38350 3522 38534
use cut_M1M4_2x2 
transform 1 0 6822 0 1 38350
box 6822 38350 7006 38534
use cut_M1M4_2x2 
transform 1 0 7298 0 1 38350
box 7298 38350 7482 38534
use cut_M1M4_2x2 
transform 1 0 10782 0 1 38350
box 10782 38350 10966 38534
use cut_M1M4_2x2 
transform 1 0 11258 0 1 38350
box 11258 38350 11442 38534
use cut_M1M4_2x2 
transform 1 0 14742 0 1 38350
box 14742 38350 14926 38534
use cut_M1M4_2x2 
transform 1 0 15218 0 1 38350
box 15218 38350 15402 38534
use cut_M1M4_2x2 
transform 1 0 18702 0 1 38350
box 18702 38350 18886 38534
use cut_M1M2_2x1 
transform 1 0 9520 0 1 450
box 9520 450 9704 518
use cut_M1M2_2x1 
transform 1 0 9520 0 1 -1380
box 9520 -1380 9704 -1312
use cut_M1M2_2x1 
transform 1 0 12520 0 1 450
box 12520 450 12704 518
use cut_M1M2_2x1 
transform 1 0 12520 0 1 -1380
box 12520 -1380 12704 -1312
use cut_M1M2_2x1 
transform 1 0 1482 0 1 34944
box 1482 34944 1666 35012
use cut_M1M2_1x2 
transform 1 0 -2032 0 1 34882
box -2032 34882 -1964 35066
use cut_M1M4_2x1 
transform 1 0 9714 0 1 -1560
box 9714 -1560 9898 -1492
use cut_M1M4_2x1 
transform 1 0 12326 0 1 -1560
box 12326 -1560 12510 -1492
use cut_M1M3_2x1 
transform 1 0 2382 0 1 35378
box 2382 35378 2566 35446
use cut_M1M3_2x1 
transform 1 0 4722 0 1 34944
box 4722 34944 4906 35012
use cut_M1M3_2x1 
transform 1 0 6342 0 1 35378
box 6342 35378 6526 35446
use cut_M1M3_2x1 
transform 1 0 8682 0 1 34944
box 8682 34944 8866 35012
use cut_M1M3_2x1 
transform 1 0 10302 0 1 35378
box 10302 35378 10486 35446
use cut_M1M3_2x1 
transform 1 0 12642 0 1 34944
box 12642 34944 12826 35012
use cut_M1M3_2x1 
transform 1 0 14262 0 1 35378
box 14262 35378 14446 35446
use cut_M1M3_2x1 
transform 1 0 16602 0 1 34944
box 16602 34944 16786 35012
use cut_M1M3_2x1 
transform 1 0 1482 0 1 32064
box 1482 32064 1666 32132
use cut_M1M3_2x1 
transform 1 0 4722 0 1 32064
box 4722 32064 4906 32132
use cut_M1M3_2x1 
transform 1 0 5442 0 1 32064
box 5442 32064 5626 32132
use cut_M1M3_2x1 
transform 1 0 8682 0 1 32064
box 8682 32064 8866 32132
use cut_M1M3_2x1 
transform 1 0 9402 0 1 32064
box 9402 32064 9586 32132
use cut_M1M3_2x1 
transform 1 0 12642 0 1 32064
box 12642 32064 12826 32132
use cut_M1M3_2x1 
transform 1 0 13362 0 1 32064
box 13362 32064 13546 32132
use cut_M1M3_2x1 
transform 1 0 16602 0 1 32064
box 16602 32064 16786 32132
use cut_M1M3_2x1 
transform 1 0 17322 0 1 32064
box 17322 32064 17506 32132
use cut_M1M2_2x1 
transform 1 0 3822 0 1 35344
box 3822 35344 4006 35412
use cut_M1M2_2x1 
transform 1 0 5442 0 1 34944
box 5442 34944 5626 35012
use cut_M1M2_2x1 
transform 1 0 7782 0 1 35344
box 7782 35344 7966 35412
use cut_M1M2_2x1 
transform 1 0 9402 0 1 34944
box 9402 34944 9586 35012
use cut_M1M2_2x1 
transform 1 0 11742 0 1 35344
box 11742 35344 11926 35412
use cut_M1M2_2x1 
transform 1 0 13362 0 1 34944
box 13362 34944 13546 35012
use cut_M1M2_2x1 
transform 1 0 15702 0 1 35344
box 15702 35344 15886 35412
use cut_M1M2_2x1 
transform 1 0 17322 0 1 34944
box 17322 34944 17506 35012
use cut_M1M3_2x1 
transform 1 0 1482 0 1 25664
box 1482 25664 1666 25732
use cut_M1M3_2x1 
transform 1 0 4722 0 1 25664
box 4722 25664 4906 25732
use cut_M1M3_2x1 
transform 1 0 5442 0 1 25664
box 5442 25664 5626 25732
use cut_M1M3_2x1 
transform 1 0 8682 0 1 25664
box 8682 25664 8866 25732
use cut_M1M3_2x1 
transform 1 0 9402 0 1 25664
box 9402 25664 9586 25732
use cut_M1M3_2x1 
transform 1 0 12642 0 1 25664
box 12642 25664 12826 25732
use cut_M1M3_2x1 
transform 1 0 13362 0 1 25664
box 13362 25664 13546 25732
use cut_M1M3_2x1 
transform 1 0 16602 0 1 25664
box 16602 25664 16786 25732
use cut_M1M3_2x1 
transform 1 0 17322 0 1 25664
box 17322 25664 17506 25732
use cut_M1M3_2x1 
transform 1 0 2742 0 1 26304
box 2742 26304 2926 26372
use cut_M1M3_2x1 
transform 1 0 2742 0 1 26304
box 2742 26304 2926 26372
use cut_M1M3_2x1 
transform 1 0 3462 0 1 26304
box 3462 26304 3646 26372
use cut_M1M3_2x1 
transform 1 0 6702 0 1 26304
box 6702 26304 6886 26372
use cut_M1M3_2x1 
transform 1 0 7422 0 1 26304
box 7422 26304 7606 26372
use cut_M1M3_2x1 
transform 1 0 10662 0 1 26304
box 10662 26304 10846 26372
use cut_M1M3_2x1 
transform 1 0 11382 0 1 26304
box 11382 26304 11566 26372
use cut_M1M3_2x1 
transform 1 0 14622 0 1 26304
box 14622 26304 14806 26372
use cut_M1M3_2x1 
transform 1 0 15342 0 1 26304
box 15342 26304 15526 26372
use cut_M1M3_2x1 
transform 1 0 18582 0 1 26304
box 18582 26304 18766 26372
use cut_M1M3_2x1 
transform 1 0 20198 0 1 27698
box 20198 27698 20382 27766
use cut_M1M3_2x1 
transform 1 0 19658 0 1 28978
box 19658 28978 19842 29046
use cut_M1M3_2x1 
transform 1 0 19302 0 1 35584
box 19302 35584 19486 35652
use cut_M1M3_2x1 
transform 1 0 17322 0 1 32704
box 17322 32704 17506 32772
use cut_M1M3_2x1 
transform 1 0 19298 0 1 36224
box 19298 36224 19482 36292
use cut_M1M3_2x1 
transform 1 0 18218 0 1 35378
box 18218 35378 18402 35446
use cut_M1M2_2x1 
transform 1 0 19298 0 1 35904
box 19298 35904 19482 35972
use cut_M1M2_2x1 
transform 1 0 17678 0 1 33424
box 17678 33424 17862 33492
use cut_M4M5_1x2 
transform 1 0 10194 0 1 1170
box 10194 1170 10262 1354
use cut_M4M5_1x2 
transform 1 0 10194 0 1 4846
box 10194 4846 10262 5030
use cut_M1M4_2x1 
transform 1 0 11742 0 1 1170
box 11742 1170 11926 1238
use cut_M4M5_1x2 
transform 1 0 11970 0 1 1170
box 11970 1170 12038 1354
use cut_M4M5_1x2 
transform 1 0 11970 0 1 4846
box 11970 4846 12038 5030
use cut_M1M3_2x1 
transform 1 0 10302 0 1 2450
box 10302 2450 10486 2518
use cut_M1M3_2x1 
transform 1 0 11742 0 1 1170
box 11742 1170 11926 1238
use cut_M1M4_2x1 
transform 1 0 10302 0 1 1170
box 10302 1170 10486 1238
use cut_M1M4_2x1 
transform 1 0 11742 0 1 2450
box 11742 2450 11926 2518
use cut_M1M3_2x1 
transform 1 0 1482 0 1 26304
box 1482 26304 1666 26372
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 5030
box -1248 5030 -1064 5214
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 6518
box -1248 6518 -1064 6702
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 8006
box -1248 8006 -1064 8190
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 9494
box -1248 9494 -1064 9678
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 10982
box -1248 10982 -1064 11166
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 12470
box -1248 12470 -1064 12654
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 13958
box -1248 13958 -1064 14142
use cut_M1M2_2x2 
transform 1 0 -1248 0 1 15446
box -1248 15446 -1064 15630
use cut_M1M2_2x2 
transform 1 0 23288 0 1 4970
box 23288 4970 23472 5154
use cut_M1M2_2x2 
transform 1 0 23288 0 1 6458
box 23288 6458 23472 6642
use cut_M1M2_2x2 
transform 1 0 23288 0 1 7946
box 23288 7946 23472 8130
use cut_M1M2_2x2 
transform 1 0 23288 0 1 9434
box 23288 9434 23472 9618
use cut_M1M2_2x2 
transform 1 0 23288 0 1 10922
box 23288 10922 23472 11106
use cut_M1M2_2x2 
transform 1 0 23288 0 1 12410
box 23288 12410 23472 12594
use cut_M1M2_2x2 
transform 1 0 23288 0 1 13898
box 23288 13898 23472 14082
use cut_M1M2_2x2 
transform 1 0 23288 0 1 15386
box 23288 15386 23472 15570
<< labels >>
flabel m3 s 1478 18634 1538 27900 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 12078 18804 12138 27922 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 16038 18974 16098 27922 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 10078 19144 10138 27922 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 14038 19314 14098 27922 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 6118 19654 6178 27922 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 4158 19824 4218 27922 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8118 19994 8178 27922 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel locali s 23288 -600 23472 37334 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
flabel locali s 23888 -1200 24072 37934 0 FreeSans 400 0 0 0 AVDD
port 10 nsew
flabel locali s -1848 38350 24072 38534 0 FreeSans 400 0 0 0 VREF
port 11 nsew
flabel locali s 24192 -1380 24252 38534 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 12 nsew
flabel locali s 17682 33424 17862 33484 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 10302 46 10486 114 0 FreeSans 400 0 0 0 SAR_IP
port 14 nsew
flabel m3 s 11738 46 11922 114 0 FreeSans 400 0 0 0 SAR_IN
port 15 nsew
flabel locali s 1482 32064 1662 32124 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 2742 26304 2922 26364 0 FreeSans 400 0 0 0 EN
port 17 nsew
flabel locali s 10302 2450 10482 2510 0 FreeSans 400 0 0 0 SARN
port 18 nsew
flabel locali s 10302 1170 10482 1230 0 FreeSans 400 0 0 0 SARP
port 19 nsew
flabel m3 s 17998 27922 18066 28106 0 FreeSans 400 0 0 0 D<0>
port 20 nsew
<< end >>
