magic
tech sky130A
magscale 1 2
timestamp 1659380236
<< checkpaint >>
rect 0 0 2520 2816
<< locali >>
rect 864 234 1032 294
rect 864 410 1032 470
rect 864 938 1032 998
rect 864 1114 1032 1174
rect 864 1642 1032 1702
rect 864 1818 1032 1878
rect 864 2346 1032 2406
rect 864 2522 1032 2582
rect 1032 234 1656 294
rect 1032 410 1656 470
rect 1032 938 1656 998
rect 1032 1114 1656 1174
rect 1032 1642 1656 1702
rect 1032 1818 1656 1878
rect 1032 2346 1656 2406
rect 1032 2522 1656 2582
rect 1032 234 1092 2582
rect 402 146 462 2670
rect 2058 146 2118 2670
rect 324 146 540 206
rect 756 234 972 294
rect 2412 132 2628 220
rect -108 132 108 220
<< poly >>
rect 324 158 2196 194
rect 324 510 2196 546
rect 324 862 2196 898
rect 324 1214 2196 1250
rect 324 1566 2196 1602
rect 324 1918 2196 1954
rect 324 2270 2196 2306
rect 324 2622 2196 2658
<< m3 >>
rect 1548 0 1748 2816
rect 756 0 956 2816
rect 1548 0 1748 2816
rect 756 0 956 2816
use SUNTRB_NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTRB_NCHDL MN1
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTRB_NCHDL MN2
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNTRB_NCHDL MN3
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNTRB_NCHDL MN4
transform 1 0 0 0 1 1408
box 0 1408 1260 1760
use SUNTRB_NCHDL MN5
transform 1 0 0 0 1 1760
box 0 1760 1260 2112
use SUNTRB_NCHDL MN6
transform 1 0 0 0 1 2112
box 0 2112 1260 2464
use SUNTRB_NCHDL MN7
transform 1 0 0 0 1 2464
box 0 2464 1260 2816
use SUNTRB_PCHDL MP0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTRB_PCHDL MP1
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTRB_PCHDL MP2
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNTRB_PCHDL MP3
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNTRB_PCHDL MP4
transform 1 0 1260 0 1 1408
box 1260 1408 2520 1760
use SUNTRB_PCHDL MP5
transform 1 0 1260 0 1 1760
box 1260 1760 2520 2112
use SUNTRB_PCHDL MP6
transform 1 0 1260 0 1 2112
box 1260 2112 2520 2464
use SUNTRB_PCHDL MP7
transform 1 0 1260 0 1 2464
box 1260 2464 2520 2816
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 586
box 1548 586 1748 662
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 762
box 1548 762 1748 838
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 1290
box 1548 1290 1748 1366
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 1466
box 1548 1466 1748 1542
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 1994
box 1548 1994 1748 2070
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 2170
box 1548 2170 1748 2246
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 2698
box 1548 2698 1748 2774
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 58
box 756 58 956 134
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 586
box 756 586 956 662
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 762
box 756 762 956 838
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 1290
box 756 1290 956 1366
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 1466
box 756 1466 956 1542
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 1994
box 756 1994 956 2070
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 2170
box 756 2170 956 2246
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 2698
box 756 2698 956 2774
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 756 234 972 294 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 3 nsew
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 4 nsew
flabel m3 s 1548 0 1748 2816 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 756 0 956 2816 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
