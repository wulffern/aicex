magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 2592 1584
<< locali >>
rect -108 -44 108 44
rect 2412 -44 2628 44
rect -108 44 108 132
rect 2412 44 2628 132
rect -108 132 108 220
rect 1692 132 1980 220
rect 1692 132 1980 220
rect 2412 132 2628 220
rect -108 220 108 308
rect 1908 220 1980 308
rect 2412 220 2628 308
rect -108 308 108 396
rect 324 308 1836 396
rect 1908 308 2196 396
rect 2412 308 2628 396
rect -108 396 108 484
rect 324 396 396 484
rect 2124 396 2196 484
rect 2412 396 2628 484
rect -108 484 108 572
rect 324 484 396 572
rect 468 484 612 572
rect 684 484 2196 572
rect 2412 484 2628 572
rect -108 572 108 660
rect 324 572 396 660
rect 2124 572 2196 660
rect 2412 572 2628 660
rect -108 660 108 748
rect 324 660 2052 748
rect 2124 660 2196 748
rect 2412 660 2628 748
rect -108 748 108 836
rect 324 748 396 836
rect 2124 748 2196 836
rect 2412 748 2628 836
rect -108 836 108 924
rect 324 836 396 924
rect 468 836 2196 924
rect 2412 836 2628 924
rect -108 924 108 1012
rect 324 924 396 1012
rect 2124 924 2196 1012
rect 2412 924 2628 1012
rect -108 1012 108 1100
rect 324 1012 1764 1100
rect 1836 1012 2052 1100
rect 2124 1012 2196 1100
rect 2412 1012 2628 1100
rect -108 1100 108 1188
rect 324 1100 396 1188
rect 2124 1100 2196 1188
rect 2412 1100 2628 1188
rect -108 1188 108 1276
rect 324 1188 828 1276
rect 900 1188 2196 1276
rect 2412 1188 2628 1276
rect -108 1276 108 1364
rect 756 1276 828 1364
rect 2412 1276 2628 1364
rect -108 1364 108 1452
rect 756 1364 2052 1452
rect 756 1364 2052 1452
rect 2412 1364 2628 1452
rect -108 1452 108 1540
rect 2412 1452 2628 1540
rect -108 1540 108 1628
rect 2412 1540 2628 1628
<< rlocali >>
rect 612 484 684 572
rect 1764 1012 1836 1100
<< labels >>
flabel locali s 1692 132 1980 220 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 756 1364 2052 1452 0 FreeSans 400 0 0 0 A
port 1 nsew
<< end >>
