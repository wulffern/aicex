magic
tech sky130A
magscale 1 2
timestamp 1658874400
<< checkpaint >>
rect 0 0 2520 5280
<< locali >>
rect 1656 586 1824 646
rect 1824 1142 2040 1202
rect 1824 586 1884 1202
rect 1980 1202 2088 1262
rect 1656 1290 1824 1350
rect 1824 1906 2088 1966
rect 1824 4722 2088 4782
rect 1824 1290 1884 4782
rect 432 2610 600 2670
rect 600 1290 864 1350
rect 600 1290 660 2670
rect 480 3606 600 3666
rect 600 1290 864 1350
rect 600 1290 660 3666
rect 432 3666 540 3726
rect 864 1994 1032 2054
rect 864 2698 1032 2758
rect 1032 1994 1092 2758
rect 432 5074 600 5134
rect 600 4810 864 4870
rect 600 4810 660 5134
rect 324 1554 540 1614
rect 324 498 540 558
rect 756 5162 972 5222
rect 756 4810 972 4870
rect 324 4018 540 4078
<< m1 >>
rect 2088 2610 2256 2670
rect 2088 3666 2256 3726
rect 1656 586 2256 646
rect 2256 586 2316 3734
rect 480 1846 600 1906
rect 600 938 864 998
rect 600 938 660 1974
rect 432 1906 540 1966
rect 864 3754 1032 3814
rect 864 4810 1032 4870
rect 1032 3754 1092 4878
rect 432 2962 600 3022
rect 600 2698 864 2758
rect 600 2698 660 3030
rect 1656 3050 1824 3110
rect 1824 2258 2088 2318
rect 1824 3314 2088 3374
rect 1824 2258 1884 3382
rect 1656 5162 1824 5222
rect 1824 4370 2088 4430
rect 1824 4370 1884 5230
rect 204 850 432 910
rect 204 4018 432 4078
rect 204 850 264 4086
<< m2 >>
rect 432 4722 604 4798
rect 604 3666 2088 3742
rect 604 3666 680 4798
<< m3 >>
rect 1548 0 1748 5280
rect 756 0 956 5280
rect 1548 0 1748 5280
rect 756 0 956 5280
use SUNTR_TAPCELLB_CV XA0
transform 1 0 0 0 1 0
box 0 0 2520 352
use SUNTR_NDX1_CV XA1
transform 1 0 0 0 1 352
box 0 352 2520 1056
use SUNTR_IVX1_CV XA2
transform 1 0 0 0 1 1056
box 0 1056 2520 1408
use SUNTR_IVTRIX1_CV XA3
transform 1 0 0 0 1 1408
box 0 1408 2520 2112
use SUNTR_IVTRIX1_CV XA4
transform 1 0 0 0 1 2112
box 0 2112 2520 2816
use SUNTR_IVX1_CV XA5
transform 1 0 0 0 1 2816
box 0 2816 2520 3168
use SUNTR_IVTRIX1_CV XA6
transform 1 0 0 0 1 3168
box 0 3168 2520 3872
use SUNTR_NDTRIX1_CV XA7
transform 1 0 0 0 1 3872
box 0 3872 2520 4928
use SUNTR_IVX1_CV XA8
transform 1 0 0 0 1 4928
box 0 4928 2520 5280
use SUNTR_cut_M1M2_2x1 
transform 1 0 1980 0 1 2610
box 1980 2610 2164 2678
use SUNTR_cut_M1M2_2x1 
transform 1 0 1980 0 1 3666
box 1980 3666 2164 3734
use SUNTR_cut_M1M2_2x1 
transform 1 0 1548 0 1 586
box 1548 586 1732 654
use SUNTR_cut_M1M2_2x1 
transform 1 0 324 0 1 1906
box 324 1906 508 1974
use SUNTR_cut_M1M2_2x1 
transform 1 0 756 0 1 938
box 756 938 940 1006
use SUNTR_cut_M1M3_2x1 
transform 1 0 324 0 1 4722
box 324 4722 524 4798
use SUNTR_cut_M1M3_2x1 
transform 1 0 1980 0 1 3666
box 1980 3666 2180 3742
use SUNTR_cut_M1M2_2x1 
transform 1 0 756 0 1 3754
box 756 3754 940 3822
use SUNTR_cut_M1M2_2x1 
transform 1 0 756 0 1 4810
box 756 4810 940 4878
use SUNTR_cut_M1M2_2x1 
transform 1 0 324 0 1 2962
box 324 2962 508 3030
use SUNTR_cut_M1M2_2x1 
transform 1 0 756 0 1 2698
box 756 2698 940 2766
use SUNTR_cut_M1M2_2x1 
transform 1 0 1548 0 1 3050
box 1548 3050 1732 3118
use SUNTR_cut_M1M2_2x1 
transform 1 0 1980 0 1 2258
box 1980 2258 2164 2326
use SUNTR_cut_M1M2_2x1 
transform 1 0 1980 0 1 3314
box 1980 3314 2164 3382
use SUNTR_cut_M1M2_2x1 
transform 1 0 1548 0 1 5162
box 1548 5162 1732 5230
use SUNTR_cut_M1M2_2x1 
transform 1 0 1980 0 1 4370
box 1980 4370 2164 4438
use SUNTR_cut_M1M2_2x1 
transform 1 0 324 0 1 850
box 324 850 508 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 324 0 1 4018
box 324 4018 508 4086
<< labels >>
flabel locali s 324 1554 540 1614 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 CK
port 2 nsew
flabel locali s 756 5162 972 5222 0 FreeSans 400 0 0 0 Q
port 4 nsew
flabel locali s 756 4810 972 4870 0 FreeSans 400 0 0 0 QN
port 5 nsew
flabel locali s 324 4018 540 4078 0 FreeSans 400 0 0 0 RN
port 3 nsew
flabel m3 s 1548 0 1748 5280 0 FreeSans 400 0 0 0 AVDD
port 6 nsew
flabel m3 s 756 0 956 5280 0 FreeSans 400 0 0 0 AVSS
port 7 nsew
<< end >>
