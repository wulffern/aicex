
*-------------------------------------------------------------
* SUNTR_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLCM D G S B
XM0 N0 G S B SUNTR_NCHDL
XM1 N1 G N0 B SUNTR_NCHDL
XM2 N2 G N1 B SUNTR_NCHDL
XM3 N3 G N2 B SUNTR_NCHDL
XM4 N4 G N3 B SUNTR_NCHDL
XM5 N5 G N4 B SUNTR_NCHDL
XM6 N6 G N5 B SUNTR_NCHDL
XM7 N7 G N6 B SUNTR_NCHDL
XM8 D G N7 B SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLCM D G S B
XM0 N0 G S B SUNTR_PCHDL
XM7 D G N0 B SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLA D G S B
XM0 D G S B SUNTR_NCHDL
XM1 S G D B SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLA D G S B
XM0 D G S B SUNTR_PCHDL
XM1 S G D B SUNTR_PCHDL
XM2 D G S B SUNTR_PCHDL
XM3 S G D B SUNTR_PCHDL
XM4 D G S B SUNTR_PCHDL
XM5 S G D B SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_RES100 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RES100 N P B
XRR1_0 N INT_0 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_1 INT_0 INT_1 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_2 INT_1 INT_2 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_3 INT_2 INT_3 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_4 INT_3 INT_4 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_5 INT_4 INT_5 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_6 INT_5 INT_6 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_7 INT_6 INT_7 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_8 INT_7 INT_8 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_9 INT_8 P B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
.ENDS

*-------------------------------------------------------------
* SUNTR_RPPO_100k <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RPPO_100k P N B
XA1 N P B SUNTR_RES100
.ENDS

*-------------------------------------------------------------
* SUNTR_TAPCELLB_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTR_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX1_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX8_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMN4 Y A AVSS AVSS SUNTR_NCHDL
XMN5 AVSS A Y AVSS SUNTR_NCHDL
XMN6 Y A AVSS AVSS SUNTR_NCHDL
XMN7 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
XMP2 Y A AVDD AVDD SUNTR_PCHDL
XMP3 AVDD A Y AVDD SUNTR_PCHDL
XMP4 Y A AVDD AVDD SUNTR_PCHDL
XMP5 AVDD A Y AVDD SUNTR_PCHDL
XMP6 Y A AVDD AVDD SUNTR_PCHDL
XMP7 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NRX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NRX1_CV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS B Y AVSS SUNTR_NCHDL
XMP0 N1 A AVDD AVDD SUNTR_PCHDL
XMP1 Y B N1 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NDX1_CV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y B N1 AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD B Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_DFTSPCX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFTSPCX1_CV D CK Q AVDD AVSS
XMN0 N1 D AVSS AVSS SUNTR_NCHDL
XMN2 N2 CK Q AVSS SUNTR_NCHDL
XMN1 AVSS N1 N2 AVSS SUNTR_NCHDL
XMP1 N3 D AVDD AVDD SUNTR_PCHDL
XMP0 N1 CK N3 AVDD SUNTR_PCHDL
XMP2 Q N1 AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVTRIX1_CV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y C N1 AVSS SUNTR_NCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NDTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NDTRIX1_CV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS SUNTR_NCHDL
XMN0 N2 A N1 AVSS SUNTR_NCHDL
XMN1 Y C N2 AVSS SUNTR_NCHDL
XMP2 AVDD RN N2 AVDD SUNTR_PCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_DFRNQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS SUNTR_TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS SUNTR_NDX1_CV
XA2 CKN CKB AVDD AVSS SUNTR_IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS SUNTR_IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS SUNTR_IVTRIX1_CV
XA5 A0 A1 AVDD AVSS SUNTR_IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS SUNTR_IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS SUNTR_NDTRIX1_CV
XA8 QN Q AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTRB_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTRB_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_IVX1_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NDX1_CV A B Y BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNTRB_NCHDL
XMN1 Y B N1 BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
XMP1 AVDD B Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_TAPCELLBAVSS_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_TAPCELLBAVSS_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTRB_NCHDL
XMP1 NC1 NC1 NC1 AVDD SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNSAR_CAP_BSSW_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNSAR_CAP_BSSW_CV A B
C1 A B 100f
.ENDS

*-------------------------------------------------------------
* CAP_LPF <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT CAP_LPF A B
C1 A B 78f
.ENDS

*-------------------------------------------------------------
* SUN_PLL_BIAS <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_BIAS IBPSR_1U PWRUP_1V8_N AVSS
xa20 IBPSR_1U PWRUP_1V8_N AVSS AVSS SUNTR_NCHDL
xa30 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa31 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa32 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa33 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa34 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa35 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa36 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa37 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa38 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
xa39 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
.ENDS

*-------------------------------------------------------------
* SUN_PLL_BUF <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_BUF AVDD VFB VI VO VBN AVSS
xa10 VS VBN AVSS AVSS SUNTR_NCHDLCM
xa20 VDP VFB VS AVSS SUNTR_NCHDLA
xa40 VGP VI VS AVSS SUNTR_NCHDLA
xc10 VGP VDP AVDD AVDD SUNTR_PCHDLA
xc20 VDP VDP AVDD AVDD SUNTR_PCHDLA
xc3_00 VO VGP AVDD AVDD SUNTR_PCHDLA
xc3_10 VO VGP AVDD AVDD SUNTR_PCHDLA
xc3_20 VO VGP AVDD AVDD SUNTR_PCHDLA
xd20 VO AVSS SUNSAR_CAP_BSSW_CV
xd30 VO AVSS SUNSAR_CAP_BSSW_CV
xd31 VO AVSS SUNSAR_CAP_BSSW_CV
xd32 VO AVSS SUNSAR_CAP_BSSW_CV
xd33 VO AVSS SUNSAR_CAP_BSSW_CV
xd34 VO AVSS SUNSAR_CAP_BSSW_CV
xd35 VO AVSS SUNSAR_CAP_BSSW_CV
xd36 VO AVSS SUNSAR_CAP_BSSW_CV
xd37 VO AVSS SUNSAR_CAP_BSSW_CV
.ENDS

*-------------------------------------------------------------
* SUN_PLL_CP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_CP AVDD CP_UP_N LPF CP_DOWN VBN AVSS LPFZ PWRUP_1V8 KICK
xa10 VBP VBN AVSS AVSS SUNTR_NCHDLCM
xa20 VNS VBN AVSS AVSS SUNTR_NCHDLCM
xa30 LPF CP_DOWN VNS AVSS SUNTR_NCHDL
xa40 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa41 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa42 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa43 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa44 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa45 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa46 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa47 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa48 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xa49 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xb10 VBP VBP AVDD AVDD SUNTR_PCHDLCM
xb20 VPS VBP AVDD AVDD SUNTR_PCHDLCM
xb30 LPF CP_UP_N VPS AVDD SUNTR_PCHDL
xb40 LPF PWRUP_1V8 AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUN_PLL_DIVN <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_DIVN AVDD CK_FB CK PWRUP_1V8 AVSS
xc0 N2 D2 PWRUP_1V8 CK_FB N2 AVDD AVSS SUNTR_DFRNQNX1_CV
xd0 N3 D3 PWRUP_1V8 D2 N3 AVDD AVSS SUNTR_DFRNQNX1_CV
xe0 N4 D4 PWRUP_1V8 D3 N4 AVDD AVSS SUNTR_DFRNQNX1_CV
xf0 N5 D5 PWRUP_1V8 D4 N5 AVDD AVSS SUNTR_DFRNQNX1_CV
xg0 N6 CK PWRUP_1V8 D5 N6 AVDD AVSS SUNTR_DFRNQNX1_CV
.ENDS

*-------------------------------------------------------------
* SUN_PLL_LPF <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_LPF VLPFZ AVSS VLPF
xa10 VN5 VLPF AVSS SUNTR_RPPO_100k
xa20 VN4 VN5 AVSS SUNTR_RPPO_100k
xa30 VN3 VN4 AVSS SUNTR_RPPO_100k
xa40 VN2 VN3 AVSS SUNTR_RPPO_100k
xa50 VLPFZ VN2 AVSS SUNTR_RPPO_100k
xb10 VLPF AVSS CAP_LPF
xb20 VLPF AVSS CAP_LPF
xb21 VLPF AVSS CAP_LPF
xb30 VLPFZ AVSS CAP_LPF
xb31 VLPFZ AVSS CAP_LPF
xb32 VLPFZ AVSS CAP_LPF
xb33 VLPFZ AVSS CAP_LPF
xb34 VLPFZ AVSS CAP_LPF
xb35 VLPFZ AVSS CAP_LPF
xb36 VLPFZ AVSS CAP_LPF
xb37 VLPFZ AVSS CAP_LPF
xb38 VLPFZ AVSS CAP_LPF
xb39 VLPFZ AVSS CAP_LPF
xb310 VLPFZ AVSS CAP_LPF
xb311 VLPFZ AVSS CAP_LPF
xb312 VLPFZ AVSS CAP_LPF
xb313 VLPFZ AVSS CAP_LPF
xb314 VLPFZ AVSS CAP_LPF
xb315 VLPFZ AVSS CAP_LPF
xb316 VLPFZ AVSS CAP_LPF
xb317 VLPFZ AVSS CAP_LPF
xb318 VLPFZ AVSS CAP_LPF
xb319 VLPFZ AVSS CAP_LPF
xb320 VLPFZ AVSS CAP_LPF
xb321 VLPFZ AVSS CAP_LPF
xb322 VLPFZ AVSS CAP_LPF
xb323 VLPFZ AVSS CAP_LPF
.ENDS

*-------------------------------------------------------------
* SUN_PLL_LSCORE <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_LSCORE A AN YN Y AVDD AVSS
xb1_00 Y AN AVSS AVSS SUNTR_NCHDL
xb1_10 Y AN AVSS AVSS SUNTR_NCHDL
xb2_00 YN A AVSS AVSS SUNTR_NCHDL
xb2_10 YN A AVSS AVSS SUNTR_NCHDL
xc1a0 net2 YN AVDD AVDD SUNTR_PCHDL
xc1b0 Y YN net2 AVDD SUNTR_PCHDL
xc2a0 net1 Y AVDD AVDD SUNTR_PCHDL
xc2b0 YN Y net1 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUN_PLL_KICK <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_KICK AVDD KICK KICK_N PWRUP_1V8 AVSS PWRUP_1V8_N
xa1a0 AVDD AVSS SUNTR_TAPCELLB_CV
xa1b0 PWRUP_1V8 PWRUP_1V8_N AVDD AVSS SUNTR_IVX1_CV
xa1c0 PWRUP_1V8_N N1 AVDD AVSS SUNTR_IVX1_CV
xa1d0 N1 __UNCONNECTED_PIN__1 AVDD AVSS SUNTR_IVX8_CV
xa20 N1 N2 AVDD AVSS SUNTR_IVX1_CV
xa3a0 N2 N3 AVDD AVSS SUNTR_IVX1_CV
xa3b0 N3 __UNCONNECTED_PIN__2 AVDD AVSS SUNTR_IVX8_CV
xa40 N3 N4 AVDD AVSS SUNTR_IVX1_CV
xa5a0 N4 N5 AVDD AVSS SUNTR_IVX1_CV
xa5b0 N5 __UNCONNECTED_PIN__3 AVDD AVSS SUNTR_IVX8_CV
xa60 N5 N6 AVDD AVSS SUNTR_IVX1_CV
xa70 N6 N7 AVDD AVSS SUNTR_IVX1_CV
xa80 PWRUP_1V8_N N7 KICK AVDD AVSS SUNTR_NRX1_CV
xa90 KICK KICK_N AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUN_PLL_PFD <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_PFD AVDD CP_UP_N CK_REF CP_DOWN CK_FB AVSS
xa00 AVDD AVSS SUNTR_TAPCELLB_CV
xa10 CFB CK_REF CP_DUP_N AVDD AVSS SUNTR_DFTSPCX1_CV
xa20 CP_DUP_N CP_UP AVDD AVSS SUNTR_IVX1_CV
xa2a0 CP_UP CP_UP_N AVDD AVSS SUNTR_IVX1_CV
xa30 CP_DUP_N CP_DOWN_N CFB AVDD AVSS SUNTR_NRX1_CV
xa50 CFB CK_FB CP_DOWN_N AVDD AVSS SUNTR_DFTSPCX1_CV
xa60 CP_DOWN_N CP_DOWN AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUN_PLL_ROSC <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_ROSC AVDD CK VDD_ROSC PWRUP_1V8 AVSS
xa3 N_2 N_1 CKUP CKDWN AVDD AVSS SUN_PLL_LSCORE
xa40 CKUP CK AVDD AVSS SUNTR_IVX1_CV
xa50 CKDWN NC1 AVDD AVSS SUNTR_IVX1_CV
xa60 AVDD AVSS SUNTR_TAPCELLB_CV
xb10 PWRUP_1V8 N_0 NI AVDD AVSS VDD_ROSC AVSS SUNTRB_NDX1_CV
xb2_00 NI N_7 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_10 N_7 N_6 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_20 N_6 N_5 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_30 N_5 N_4 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_40 N_4 N_3 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_50 N_3 N_2 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_60 N_2 N_1 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_70 N_1 N_0 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb30 AVDD AVSS SUNTRB_TAPCELLBAVSS_CV
.ENDS

*-------------------------------------------------------------
* SUN_PLL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U
xb1 AVDD VDD_ROSC VLPF VDD_ROSC IBPSR_1U AVSS SUN_PLL_BUF
xb2 VLPFZ AVSS VLPF SUN_PLL_LPF
xc1 AVDD CK_FB CK PWRUP_1V8 AVSS SUN_PLL_DIVN
xd1 AVDD CK VDD_ROSC PWRUP_1V8 AVSS SUN_PLL_ROSC
xk1 AVDD KICK __UNCONNECTED_PIN__0 PWRUP_1V8 AVSS PWRUP_1V8_N SUN_PLL_KICK
xk2 AVDD CP_UP_N VLPF CP_DOWN IBPSR_1U AVSS VLPFZ PWRUP_1V8 KICK SUN_PLL_CP
xk3 AVDD CP_UP_N CK_REF CP_DOWN CK_FB AVSS SUN_PLL_PFD
xl1 IBPSR_1U PWRUP_1V8_N AVSS SUN_PLL_BIAS
.ENDS
