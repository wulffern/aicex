magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect -600 -1080 600 1320
<< locali >>
rect -600 -1080 600 -896
rect -600 1136 600 1320
rect -600 -1080 -416 1320
rect 416 -1080 600 1320
<< labels >>
<< end >>
