magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 320
<< locali >>
rect 360 130 514 190
rect 514 210 720 270
rect 514 130 574 270
rect 1290 210 1470 270
<< poly >>
rect 270 142 1830 178
<< m3 >>
rect 1290 0 1474 320
rect 630 0 814 320
rect 1290 0 1474 320
rect 630 0 814 320
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use cut_M1M4_2x1 
transform 1 0 1290 0 1 50
box 1290 50 1474 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
<< labels >>
flabel locali s 1290 210 1470 270 0 FreeSans 400 0 0 0 Y
port 1 nsew
flabel m3 s 1290 0 1474 320 0 FreeSans 400 0 0 0 AVDD
port 2 nsew
flabel m3 s 630 0 814 320 0 FreeSans 400 0 0 0 AVSS
port 3 nsew
<< end >>
