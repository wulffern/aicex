magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 5384 4140
<< locali >>
rect 0 0 5384 112
rect 0 0 5384 112
rect 0 0 112 4140
rect 0 4028 5384 4140
rect 5272 0 5384 4140
rect 0 0 5384 112
rect 4474 3390 4798 3610
rect 586 3390 910 3610
<< ptapc >>
rect 12 0 92 80
rect 92 0 172 80
rect 172 0 252 80
rect 252 0 332 80
rect 332 0 412 80
rect 412 0 492 80
rect 492 0 572 80
rect 572 0 652 80
rect 652 0 732 80
rect 732 0 812 80
rect 812 0 892 80
rect 892 0 972 80
rect 972 0 1052 80
rect 1052 0 1132 80
rect 1132 0 1212 80
rect 1212 0 1292 80
rect 1292 0 1372 80
rect 1372 0 1452 80
rect 1452 0 1532 80
rect 1532 0 1612 80
rect 1612 0 1692 80
rect 1692 0 1772 80
rect 1772 0 1852 80
rect 1852 0 1932 80
rect 1932 0 2012 80
rect 2012 0 2092 80
rect 2092 0 2172 80
rect 2172 0 2252 80
rect 2252 0 2332 80
rect 2332 0 2412 80
rect 2412 0 2492 80
rect 2492 0 2572 80
rect 2572 0 2652 80
rect 2652 0 2732 80
rect 2732 0 2812 80
rect 2812 0 2892 80
rect 2892 0 2972 80
rect 2972 0 3052 80
rect 3052 0 3132 80
rect 3132 0 3212 80
rect 3212 0 3292 80
rect 3292 0 3372 80
rect 3372 0 3452 80
rect 3452 0 3532 80
rect 3532 0 3612 80
rect 3612 0 3692 80
rect 3692 0 3772 80
rect 3772 0 3852 80
rect 3852 0 3932 80
rect 3932 0 4012 80
rect 4012 0 4092 80
rect 4092 0 4172 80
rect 4172 0 4252 80
rect 4252 0 4332 80
rect 4332 0 4412 80
rect 4412 0 4492 80
rect 4492 0 4572 80
rect 4572 0 4652 80
rect 4652 0 4732 80
rect 4732 0 4812 80
rect 4812 0 4892 80
rect 4892 0 4972 80
rect 4972 0 5052 80
rect 5052 0 5132 80
rect 5132 0 5212 80
rect 5212 0 5292 80
rect 5292 0 5372 80
rect 0 30 80 110
rect 0 110 80 190
rect 0 190 80 270
rect 0 270 80 350
rect 0 350 80 430
rect 0 430 80 510
rect 0 510 80 590
rect 0 590 80 670
rect 0 670 80 750
rect 0 750 80 830
rect 0 830 80 910
rect 0 910 80 990
rect 0 990 80 1070
rect 0 1070 80 1150
rect 0 1150 80 1230
rect 0 1230 80 1310
rect 0 1310 80 1390
rect 0 1390 80 1470
rect 0 1470 80 1550
rect 0 1550 80 1630
rect 0 1630 80 1710
rect 0 1710 80 1790
rect 0 1790 80 1870
rect 0 1870 80 1950
rect 0 1950 80 2030
rect 0 2030 80 2110
rect 0 2110 80 2190
rect 0 2190 80 2270
rect 0 2270 80 2350
rect 0 2350 80 2430
rect 0 2430 80 2510
rect 0 2510 80 2590
rect 0 2590 80 2670
rect 0 2670 80 2750
rect 0 2750 80 2830
rect 0 2830 80 2910
rect 0 2910 80 2990
rect 0 2990 80 3070
rect 0 3070 80 3150
rect 0 3150 80 3230
rect 0 3230 80 3310
rect 0 3310 80 3390
rect 0 3390 80 3470
rect 0 3470 80 3550
rect 0 3550 80 3630
rect 0 3630 80 3710
rect 0 3710 80 3790
rect 0 3790 80 3870
rect 0 3870 80 3950
rect 0 3950 80 4030
rect 0 4030 80 4110
rect 12 4028 92 4108
rect 92 4028 172 4108
rect 172 4028 252 4108
rect 252 4028 332 4108
rect 332 4028 412 4108
rect 412 4028 492 4108
rect 492 4028 572 4108
rect 572 4028 652 4108
rect 652 4028 732 4108
rect 732 4028 812 4108
rect 812 4028 892 4108
rect 892 4028 972 4108
rect 972 4028 1052 4108
rect 1052 4028 1132 4108
rect 1132 4028 1212 4108
rect 1212 4028 1292 4108
rect 1292 4028 1372 4108
rect 1372 4028 1452 4108
rect 1452 4028 1532 4108
rect 1532 4028 1612 4108
rect 1612 4028 1692 4108
rect 1692 4028 1772 4108
rect 1772 4028 1852 4108
rect 1852 4028 1932 4108
rect 1932 4028 2012 4108
rect 2012 4028 2092 4108
rect 2092 4028 2172 4108
rect 2172 4028 2252 4108
rect 2252 4028 2332 4108
rect 2332 4028 2412 4108
rect 2412 4028 2492 4108
rect 2492 4028 2572 4108
rect 2572 4028 2652 4108
rect 2652 4028 2732 4108
rect 2732 4028 2812 4108
rect 2812 4028 2892 4108
rect 2892 4028 2972 4108
rect 2972 4028 3052 4108
rect 3052 4028 3132 4108
rect 3132 4028 3212 4108
rect 3212 4028 3292 4108
rect 3292 4028 3372 4108
rect 3372 4028 3452 4108
rect 3452 4028 3532 4108
rect 3532 4028 3612 4108
rect 3612 4028 3692 4108
rect 3692 4028 3772 4108
rect 3772 4028 3852 4108
rect 3852 4028 3932 4108
rect 3932 4028 4012 4108
rect 4012 4028 4092 4108
rect 4092 4028 4172 4108
rect 4172 4028 4252 4108
rect 4252 4028 4332 4108
rect 4332 4028 4412 4108
rect 4412 4028 4492 4108
rect 4492 4028 4572 4108
rect 4572 4028 4652 4108
rect 4652 4028 4732 4108
rect 4732 4028 4812 4108
rect 4812 4028 4892 4108
rect 4892 4028 4972 4108
rect 4972 4028 5052 4108
rect 5052 4028 5132 4108
rect 5132 4028 5212 4108
rect 5212 4028 5292 4108
rect 5292 4028 5372 4108
rect 5272 30 5352 110
rect 5272 110 5352 190
rect 5272 190 5352 270
rect 5272 270 5352 350
rect 5272 350 5352 430
rect 5272 430 5352 510
rect 5272 510 5352 590
rect 5272 590 5352 670
rect 5272 670 5352 750
rect 5272 750 5352 830
rect 5272 830 5352 910
rect 5272 910 5352 990
rect 5272 990 5352 1070
rect 5272 1070 5352 1150
rect 5272 1150 5352 1230
rect 5272 1230 5352 1310
rect 5272 1310 5352 1390
rect 5272 1390 5352 1470
rect 5272 1470 5352 1550
rect 5272 1550 5352 1630
rect 5272 1630 5352 1710
rect 5272 1710 5352 1790
rect 5272 1790 5352 1870
rect 5272 1870 5352 1950
rect 5272 1950 5352 2030
rect 5272 2030 5352 2110
rect 5272 2110 5352 2190
rect 5272 2190 5352 2270
rect 5272 2270 5352 2350
rect 5272 2350 5352 2430
rect 5272 2430 5352 2510
rect 5272 2510 5352 2590
rect 5272 2590 5352 2670
rect 5272 2670 5352 2750
rect 5272 2750 5352 2830
rect 5272 2830 5352 2910
rect 5272 2910 5352 2990
rect 5272 2990 5352 3070
rect 5272 3070 5352 3150
rect 5272 3150 5352 3230
rect 5272 3230 5352 3310
rect 5272 3310 5352 3390
rect 5272 3390 5352 3470
rect 5272 3470 5352 3550
rect 5272 3550 5352 3630
rect 5272 3630 5352 3710
rect 5272 3710 5352 3790
rect 5272 3790 5352 3870
rect 5272 3870 5352 3950
rect 5272 3950 5352 4030
rect 5272 4030 5352 4110
<< ptap >>
rect 0 0 5384 112
rect 0 0 112 4140
rect 0 4028 5384 4140
rect 5272 0 5384 4140
use SUNTR_RES200 XA1
transform 1 0 640 0 1 640
box 640 640 4744 3500
<< labels >>
flabel locali s 0 0 5384 112 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 4474 3390 4798 3610 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 586 3390 910 3610 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
