magic
tech sky130A
magscale 1 2
timestamp 1658699483
<< checkpaint >>
rect 112 0 11844 22780
<< m1 >>
rect 2100 8660 2160 22720
rect 2100 8660 2160 22720
rect 1920 140 1980 22720
rect 1920 140 1980 22720
rect 1740 17180 1800 22720
rect 1740 17180 1800 22720
rect 1560 2980 1620 22720
rect 1560 2980 1620 22720
rect 1380 6304 1440 22720
rect 1380 6304 1440 22720
rect 1200 14824 1260 22720
rect 1200 14824 1260 22720
rect 1020 14340 1080 22720
rect 1020 14340 1080 22720
rect 840 15792 900 22720
rect 840 15792 900 22720
rect 660 7272 720 22720
rect 660 7272 720 22720
rect 480 7756 540 22720
rect 480 7756 540 22720
rect 300 6788 360 22720
rect 300 6788 360 22720
rect 120 8240 180 22720
rect 120 8240 180 22720
rect 2668 0 11768 76
<< m2 >>
rect 2160 8722 2340 8798
rect 2160 11142 2340 11218
rect 2160 9690 2340 9766
rect 2160 10658 2340 10734
rect 2160 10174 2340 10250
rect 2160 9206 2340 9282
rect 2160 8722 2340 8798
rect 2160 11142 2340 11218
rect 2160 9690 2340 9766
rect 2160 10658 2340 10734
rect 2160 10174 2340 10250
rect 2160 9206 2340 9282
rect 2160 8722 2340 8798
rect 2160 11142 2340 11218
rect 2160 9690 2340 9766
rect 2160 10658 2340 10734
rect 2160 10174 2340 10250
rect 2160 9206 2340 9282
rect 2160 8722 2340 8798
rect 2160 11142 2340 11218
rect 2160 9690 2340 9766
rect 2160 10658 2340 10734
rect 2160 10174 2340 10250
rect 2160 9206 2340 9282
rect 2160 8722 2340 8798
rect 2160 11142 2340 11218
rect 2160 9690 2340 9766
rect 2160 10658 2340 10734
rect 2160 10174 2340 10250
rect 2160 9206 2340 9282
rect 2160 8722 2340 8798
rect 2160 11142 2340 11218
rect 2160 9690 2340 9766
rect 2160 10658 2340 10734
rect 2160 10174 2340 10250
rect 2160 9206 2340 9282
rect 2160 20082 2340 20158
rect 2160 22502 2340 22578
rect 2160 21050 2340 21126
rect 2160 22018 2340 22094
rect 2160 21534 2340 21610
rect 2160 20566 2340 20642
rect 2160 20082 2340 20158
rect 2160 22502 2340 22578
rect 2160 21050 2340 21126
rect 2160 22018 2340 22094
rect 2160 21534 2340 21610
rect 2160 20566 2340 20642
rect 2160 20082 2340 20158
rect 2160 22502 2340 22578
rect 2160 21050 2340 21126
rect 2160 22018 2340 22094
rect 2160 21534 2340 21610
rect 2160 20566 2340 20642
rect 2160 20082 2340 20158
rect 2160 22502 2340 22578
rect 2160 21050 2340 21126
rect 2160 22018 2340 22094
rect 2160 21534 2340 21610
rect 2160 20566 2340 20642
rect 2160 20082 2340 20158
rect 2160 22502 2340 22578
rect 2160 21050 2340 21126
rect 2160 22018 2340 22094
rect 2160 21534 2340 21610
rect 2160 20566 2340 20642
rect 2160 20082 2340 20158
rect 2160 22502 2340 22578
rect 2160 21050 2340 21126
rect 2160 22018 2340 22094
rect 2160 21534 2340 21610
rect 2160 20566 2340 20642
rect 1980 202 2340 278
rect 1980 2622 2340 2698
rect 1980 1170 2340 1246
rect 1980 2138 2340 2214
rect 1980 1654 2340 1730
rect 1980 686 2340 762
rect 1980 202 2340 278
rect 1980 2622 2340 2698
rect 1980 1170 2340 1246
rect 1980 2138 2340 2214
rect 1980 1654 2340 1730
rect 1980 686 2340 762
rect 1980 202 2340 278
rect 1980 2622 2340 2698
rect 1980 1170 2340 1246
rect 1980 2138 2340 2214
rect 1980 1654 2340 1730
rect 1980 686 2340 762
rect 1980 202 2340 278
rect 1980 2622 2340 2698
rect 1980 1170 2340 1246
rect 1980 2138 2340 2214
rect 1980 1654 2340 1730
rect 1980 686 2340 762
rect 1980 202 2340 278
rect 1980 2622 2340 2698
rect 1980 1170 2340 1246
rect 1980 2138 2340 2214
rect 1980 1654 2340 1730
rect 1980 686 2340 762
rect 1980 202 2340 278
rect 1980 2622 2340 2698
rect 1980 1170 2340 1246
rect 1980 2138 2340 2214
rect 1980 1654 2340 1730
rect 1980 686 2340 762
rect 1980 11562 2340 11638
rect 1980 13982 2340 14058
rect 1980 12530 2340 12606
rect 1980 13498 2340 13574
rect 1980 13014 2340 13090
rect 1980 12046 2340 12122
rect 1980 11562 2340 11638
rect 1980 13982 2340 14058
rect 1980 12530 2340 12606
rect 1980 13498 2340 13574
rect 1980 13014 2340 13090
rect 1980 12046 2340 12122
rect 1980 11562 2340 11638
rect 1980 13982 2340 14058
rect 1980 12530 2340 12606
rect 1980 13498 2340 13574
rect 1980 13014 2340 13090
rect 1980 12046 2340 12122
rect 1980 11562 2340 11638
rect 1980 13982 2340 14058
rect 1980 12530 2340 12606
rect 1980 13498 2340 13574
rect 1980 13014 2340 13090
rect 1980 12046 2340 12122
rect 1980 11562 2340 11638
rect 1980 13982 2340 14058
rect 1980 12530 2340 12606
rect 1980 13498 2340 13574
rect 1980 13014 2340 13090
rect 1980 12046 2340 12122
rect 1980 11562 2340 11638
rect 1980 13982 2340 14058
rect 1980 12530 2340 12606
rect 1980 13498 2340 13574
rect 1980 13014 2340 13090
rect 1980 12046 2340 12122
rect 1800 17242 2340 17318
rect 1800 19662 2340 19738
rect 1800 18210 2340 18286
rect 1800 19178 2340 19254
rect 1800 18694 2340 18770
rect 1800 17726 2340 17802
rect 1800 17242 2340 17318
rect 1800 19662 2340 19738
rect 1800 18210 2340 18286
rect 1800 19178 2340 19254
rect 1800 18694 2340 18770
rect 1800 17726 2340 17802
rect 1800 17242 2340 17318
rect 1800 19662 2340 19738
rect 1800 18210 2340 18286
rect 1800 19178 2340 19254
rect 1800 18694 2340 18770
rect 1800 17726 2340 17802
rect 1800 17242 2340 17318
rect 1800 19662 2340 19738
rect 1800 18210 2340 18286
rect 1800 19178 2340 19254
rect 1800 18694 2340 18770
rect 1800 17726 2340 17802
rect 1800 17242 2340 17318
rect 1800 19662 2340 19738
rect 1800 18210 2340 18286
rect 1800 19178 2340 19254
rect 1800 18694 2340 18770
rect 1800 17726 2340 17802
rect 1800 17242 2340 17318
rect 1800 19662 2340 19738
rect 1800 18210 2340 18286
rect 1800 19178 2340 19254
rect 1800 18694 2340 18770
rect 1800 17726 2340 17802
rect 1620 3042 2340 3118
rect 1620 5462 2340 5538
rect 1620 4010 2340 4086
rect 1620 4978 2340 5054
rect 1620 4494 2340 4570
rect 1620 3526 2340 3602
rect 1620 3042 2340 3118
rect 1620 5462 2340 5538
rect 1620 4010 2340 4086
rect 1620 4978 2340 5054
rect 1620 4494 2340 4570
rect 1620 3526 2340 3602
rect 1620 3042 2340 3118
rect 1620 5462 2340 5538
rect 1620 4010 2340 4086
rect 1620 4978 2340 5054
rect 1620 4494 2340 4570
rect 1620 3526 2340 3602
rect 1620 3042 2340 3118
rect 1620 5462 2340 5538
rect 1620 4010 2340 4086
rect 1620 4978 2340 5054
rect 1620 4494 2340 4570
rect 1620 3526 2340 3602
rect 1620 3042 2340 3118
rect 1620 5462 2340 5538
rect 1620 4010 2340 4086
rect 1620 4978 2340 5054
rect 1620 4494 2340 4570
rect 1620 3526 2340 3602
rect 1620 3042 2340 3118
rect 1620 5462 2340 5538
rect 1620 4010 2340 4086
rect 1620 4978 2340 5054
rect 1620 4494 2340 4570
rect 1620 3526 2340 3602
rect 1440 6366 2340 6442
rect 1260 14886 2340 14962
rect 1080 14402 2340 14478
rect 1080 16822 2340 16898
rect 1080 15370 2340 15446
rect 1080 16338 2340 16414
rect 1080 14402 2340 14478
rect 1080 16822 2340 16898
rect 1080 15370 2340 15446
rect 1080 16338 2340 16414
rect 1080 14402 2340 14478
rect 1080 16822 2340 16898
rect 1080 15370 2340 15446
rect 1080 16338 2340 16414
rect 1080 14402 2340 14478
rect 1080 16822 2340 16898
rect 1080 15370 2340 15446
rect 1080 16338 2340 16414
rect 900 15854 2340 15930
rect 720 7334 2340 7410
rect 540 7818 2340 7894
rect 360 6850 2340 6926
rect 180 8302 2340 8378
<< m3 >>
rect 2668 19880 2744 22780
use CAP32C_CV XC1
transform 1 0 2340 0 1 0
box 2340 0 11844 2840
use CAP32C_CV XC64a<0>
transform 1 0 2340 0 1 2840
box 2340 2840 11844 5680
use CAP32C_CV XC32a<0>
transform 1 0 2340 0 1 5680
box 2340 5680 11844 8520
use CAP32C_CV XC128a<1>
transform 1 0 2340 0 1 8520
box 2340 8520 11844 11360
use CAP32C_CV XC128b<2>
transform 1 0 2340 0 1 11360
box 2340 11360 11844 14200
use CAP32C_CV X16ab
transform 1 0 2340 0 1 14200
box 2340 14200 11844 17040
use CAP32C_CV XC64b<1>
transform 1 0 2340 0 1 17040
box 2340 17040 11844 19880
use CAP32C_CV XC0
transform 1 0 2340 0 1 19880
box 2340 19880 11844 22720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8722
box 2340 8722 2540 8798
use cut_M2M3_1x2 
transform 1 0 2092 0 1 8660
box 2092 8660 2168 8860
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11142
box 2340 11142 2540 11218
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11080
box 2092 11080 2168 11280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9690
box 2340 9690 2540 9766
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9628
box 2092 9628 2168 9828
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10658
box 2340 10658 2540 10734
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10596
box 2092 10596 2168 10796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10174
box 2340 10174 2540 10250
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10112
box 2092 10112 2168 10312
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9206
box 2340 9206 2540 9282
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9144
box 2092 9144 2168 9344
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8722
box 2340 8722 2540 8798
use cut_M2M3_1x2 
transform 1 0 2092 0 1 8660
box 2092 8660 2168 8860
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11142
box 2340 11142 2540 11218
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11080
box 2092 11080 2168 11280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9690
box 2340 9690 2540 9766
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9628
box 2092 9628 2168 9828
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10658
box 2340 10658 2540 10734
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10596
box 2092 10596 2168 10796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10174
box 2340 10174 2540 10250
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10112
box 2092 10112 2168 10312
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9206
box 2340 9206 2540 9282
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9144
box 2092 9144 2168 9344
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8722
box 2340 8722 2540 8798
use cut_M2M3_1x2 
transform 1 0 2092 0 1 8660
box 2092 8660 2168 8860
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11142
box 2340 11142 2540 11218
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11080
box 2092 11080 2168 11280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9690
box 2340 9690 2540 9766
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9628
box 2092 9628 2168 9828
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10658
box 2340 10658 2540 10734
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10596
box 2092 10596 2168 10796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10174
box 2340 10174 2540 10250
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10112
box 2092 10112 2168 10312
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9206
box 2340 9206 2540 9282
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9144
box 2092 9144 2168 9344
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8722
box 2340 8722 2540 8798
use cut_M2M3_1x2 
transform 1 0 2092 0 1 8660
box 2092 8660 2168 8860
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11142
box 2340 11142 2540 11218
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11080
box 2092 11080 2168 11280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9690
box 2340 9690 2540 9766
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9628
box 2092 9628 2168 9828
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10658
box 2340 10658 2540 10734
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10596
box 2092 10596 2168 10796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10174
box 2340 10174 2540 10250
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10112
box 2092 10112 2168 10312
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9206
box 2340 9206 2540 9282
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9144
box 2092 9144 2168 9344
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8722
box 2340 8722 2540 8798
use cut_M2M3_1x2 
transform 1 0 2092 0 1 8660
box 2092 8660 2168 8860
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11142
box 2340 11142 2540 11218
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11080
box 2092 11080 2168 11280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9690
box 2340 9690 2540 9766
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9628
box 2092 9628 2168 9828
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10658
box 2340 10658 2540 10734
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10596
box 2092 10596 2168 10796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10174
box 2340 10174 2540 10250
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10112
box 2092 10112 2168 10312
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9206
box 2340 9206 2540 9282
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9144
box 2092 9144 2168 9344
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8722
box 2340 8722 2540 8798
use cut_M2M3_1x2 
transform 1 0 2092 0 1 8660
box 2092 8660 2168 8860
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11142
box 2340 11142 2540 11218
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11080
box 2092 11080 2168 11280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9690
box 2340 9690 2540 9766
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9628
box 2092 9628 2168 9828
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10658
box 2340 10658 2540 10734
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10596
box 2092 10596 2168 10796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10174
box 2340 10174 2540 10250
use cut_M2M3_1x2 
transform 1 0 2092 0 1 10112
box 2092 10112 2168 10312
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9206
box 2340 9206 2540 9282
use cut_M2M3_1x2 
transform 1 0 2092 0 1 9144
box 2092 9144 2168 9344
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20082
box 2340 20082 2540 20158
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20020
box 2092 20020 2168 20220
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22502
box 2340 22502 2540 22578
use cut_M2M3_1x2 
transform 1 0 2092 0 1 22440
box 2092 22440 2168 22640
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21050
box 2340 21050 2540 21126
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20988
box 2092 20988 2168 21188
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22018
box 2340 22018 2540 22094
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21956
box 2092 21956 2168 22156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21534
box 2340 21534 2540 21610
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21472
box 2092 21472 2168 21672
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20566
box 2340 20566 2540 20642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20504
box 2092 20504 2168 20704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20082
box 2340 20082 2540 20158
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20020
box 2092 20020 2168 20220
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22502
box 2340 22502 2540 22578
use cut_M2M3_1x2 
transform 1 0 2092 0 1 22440
box 2092 22440 2168 22640
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21050
box 2340 21050 2540 21126
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20988
box 2092 20988 2168 21188
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22018
box 2340 22018 2540 22094
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21956
box 2092 21956 2168 22156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21534
box 2340 21534 2540 21610
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21472
box 2092 21472 2168 21672
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20566
box 2340 20566 2540 20642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20504
box 2092 20504 2168 20704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20082
box 2340 20082 2540 20158
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20020
box 2092 20020 2168 20220
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22502
box 2340 22502 2540 22578
use cut_M2M3_1x2 
transform 1 0 2092 0 1 22440
box 2092 22440 2168 22640
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21050
box 2340 21050 2540 21126
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20988
box 2092 20988 2168 21188
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22018
box 2340 22018 2540 22094
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21956
box 2092 21956 2168 22156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21534
box 2340 21534 2540 21610
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21472
box 2092 21472 2168 21672
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20566
box 2340 20566 2540 20642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20504
box 2092 20504 2168 20704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20082
box 2340 20082 2540 20158
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20020
box 2092 20020 2168 20220
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22502
box 2340 22502 2540 22578
use cut_M2M3_1x2 
transform 1 0 2092 0 1 22440
box 2092 22440 2168 22640
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21050
box 2340 21050 2540 21126
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20988
box 2092 20988 2168 21188
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22018
box 2340 22018 2540 22094
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21956
box 2092 21956 2168 22156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21534
box 2340 21534 2540 21610
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21472
box 2092 21472 2168 21672
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20566
box 2340 20566 2540 20642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20504
box 2092 20504 2168 20704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20082
box 2340 20082 2540 20158
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20020
box 2092 20020 2168 20220
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22502
box 2340 22502 2540 22578
use cut_M2M3_1x2 
transform 1 0 2092 0 1 22440
box 2092 22440 2168 22640
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21050
box 2340 21050 2540 21126
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20988
box 2092 20988 2168 21188
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22018
box 2340 22018 2540 22094
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21956
box 2092 21956 2168 22156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21534
box 2340 21534 2540 21610
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21472
box 2092 21472 2168 21672
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20566
box 2340 20566 2540 20642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20504
box 2092 20504 2168 20704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20082
box 2340 20082 2540 20158
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20020
box 2092 20020 2168 20220
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22502
box 2340 22502 2540 22578
use cut_M2M3_1x2 
transform 1 0 2092 0 1 22440
box 2092 22440 2168 22640
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21050
box 2340 21050 2540 21126
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20988
box 2092 20988 2168 21188
use cut_M1M3_2x1 
transform 1 0 2340 0 1 22018
box 2340 22018 2540 22094
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21956
box 2092 21956 2168 22156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 21534
box 2340 21534 2540 21610
use cut_M2M3_1x2 
transform 1 0 2092 0 1 21472
box 2092 21472 2168 21672
use cut_M1M3_2x1 
transform 1 0 2340 0 1 20566
box 2340 20566 2540 20642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 20504
box 2092 20504 2168 20704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2622
box 2340 2622 2540 2698
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2560
box 1912 2560 1988 2760
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1170
box 2340 1170 2540 1246
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1108
box 1912 1108 1988 1308
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2138
box 2340 2138 2540 2214
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2076
box 1912 2076 1988 2276
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1654
box 2340 1654 2540 1730
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1592
box 1912 1592 1988 1792
use cut_M1M3_2x1 
transform 1 0 2340 0 1 686
box 2340 686 2540 762
use cut_M2M3_1x2 
transform 1 0 1912 0 1 624
box 1912 624 1988 824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2622
box 2340 2622 2540 2698
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2560
box 1912 2560 1988 2760
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1170
box 2340 1170 2540 1246
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1108
box 1912 1108 1988 1308
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2138
box 2340 2138 2540 2214
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2076
box 1912 2076 1988 2276
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1654
box 2340 1654 2540 1730
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1592
box 1912 1592 1988 1792
use cut_M1M3_2x1 
transform 1 0 2340 0 1 686
box 2340 686 2540 762
use cut_M2M3_1x2 
transform 1 0 1912 0 1 624
box 1912 624 1988 824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2622
box 2340 2622 2540 2698
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2560
box 1912 2560 1988 2760
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1170
box 2340 1170 2540 1246
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1108
box 1912 1108 1988 1308
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2138
box 2340 2138 2540 2214
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2076
box 1912 2076 1988 2276
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1654
box 2340 1654 2540 1730
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1592
box 1912 1592 1988 1792
use cut_M1M3_2x1 
transform 1 0 2340 0 1 686
box 2340 686 2540 762
use cut_M2M3_1x2 
transform 1 0 1912 0 1 624
box 1912 624 1988 824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2622
box 2340 2622 2540 2698
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2560
box 1912 2560 1988 2760
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1170
box 2340 1170 2540 1246
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1108
box 1912 1108 1988 1308
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2138
box 2340 2138 2540 2214
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2076
box 1912 2076 1988 2276
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1654
box 2340 1654 2540 1730
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1592
box 1912 1592 1988 1792
use cut_M1M3_2x1 
transform 1 0 2340 0 1 686
box 2340 686 2540 762
use cut_M2M3_1x2 
transform 1 0 1912 0 1 624
box 1912 624 1988 824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2622
box 2340 2622 2540 2698
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2560
box 1912 2560 1988 2760
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1170
box 2340 1170 2540 1246
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1108
box 1912 1108 1988 1308
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2138
box 2340 2138 2540 2214
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2076
box 1912 2076 1988 2276
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1654
box 2340 1654 2540 1730
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1592
box 1912 1592 1988 1792
use cut_M1M3_2x1 
transform 1 0 2340 0 1 686
box 2340 686 2540 762
use cut_M2M3_1x2 
transform 1 0 1912 0 1 624
box 1912 624 1988 824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2622
box 2340 2622 2540 2698
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2560
box 1912 2560 1988 2760
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1170
box 2340 1170 2540 1246
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1108
box 1912 1108 1988 1308
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2138
box 2340 2138 2540 2214
use cut_M2M3_1x2 
transform 1 0 1912 0 1 2076
box 1912 2076 1988 2276
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1654
box 2340 1654 2540 1730
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1592
box 1912 1592 1988 1792
use cut_M1M3_2x1 
transform 1 0 2340 0 1 686
box 2340 686 2540 762
use cut_M2M3_1x2 
transform 1 0 1912 0 1 624
box 1912 624 1988 824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11562
box 2340 11562 2540 11638
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11500
box 1912 11500 1988 11700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13982
box 2340 13982 2540 14058
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13920
box 1912 13920 1988 14120
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12530
box 2340 12530 2540 12606
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12468
box 1912 12468 1988 12668
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13498
box 2340 13498 2540 13574
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13436
box 1912 13436 1988 13636
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13014
box 2340 13014 2540 13090
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12952
box 1912 12952 1988 13152
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12046
box 2340 12046 2540 12122
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11984
box 1912 11984 1988 12184
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11562
box 2340 11562 2540 11638
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11500
box 1912 11500 1988 11700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13982
box 2340 13982 2540 14058
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13920
box 1912 13920 1988 14120
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12530
box 2340 12530 2540 12606
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12468
box 1912 12468 1988 12668
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13498
box 2340 13498 2540 13574
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13436
box 1912 13436 1988 13636
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13014
box 2340 13014 2540 13090
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12952
box 1912 12952 1988 13152
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12046
box 2340 12046 2540 12122
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11984
box 1912 11984 1988 12184
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11562
box 2340 11562 2540 11638
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11500
box 1912 11500 1988 11700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13982
box 2340 13982 2540 14058
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13920
box 1912 13920 1988 14120
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12530
box 2340 12530 2540 12606
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12468
box 1912 12468 1988 12668
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13498
box 2340 13498 2540 13574
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13436
box 1912 13436 1988 13636
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13014
box 2340 13014 2540 13090
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12952
box 1912 12952 1988 13152
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12046
box 2340 12046 2540 12122
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11984
box 1912 11984 1988 12184
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11562
box 2340 11562 2540 11638
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11500
box 1912 11500 1988 11700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13982
box 2340 13982 2540 14058
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13920
box 1912 13920 1988 14120
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12530
box 2340 12530 2540 12606
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12468
box 1912 12468 1988 12668
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13498
box 2340 13498 2540 13574
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13436
box 1912 13436 1988 13636
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13014
box 2340 13014 2540 13090
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12952
box 1912 12952 1988 13152
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12046
box 2340 12046 2540 12122
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11984
box 1912 11984 1988 12184
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11562
box 2340 11562 2540 11638
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11500
box 1912 11500 1988 11700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13982
box 2340 13982 2540 14058
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13920
box 1912 13920 1988 14120
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12530
box 2340 12530 2540 12606
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12468
box 1912 12468 1988 12668
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13498
box 2340 13498 2540 13574
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13436
box 1912 13436 1988 13636
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13014
box 2340 13014 2540 13090
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12952
box 1912 12952 1988 13152
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12046
box 2340 12046 2540 12122
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11984
box 1912 11984 1988 12184
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11562
box 2340 11562 2540 11638
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11500
box 1912 11500 1988 11700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13982
box 2340 13982 2540 14058
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13920
box 1912 13920 1988 14120
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12530
box 2340 12530 2540 12606
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12468
box 1912 12468 1988 12668
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13498
box 2340 13498 2540 13574
use cut_M2M3_1x2 
transform 1 0 1912 0 1 13436
box 1912 13436 1988 13636
use cut_M1M3_2x1 
transform 1 0 2340 0 1 13014
box 2340 13014 2540 13090
use cut_M2M3_1x2 
transform 1 0 1912 0 1 12952
box 1912 12952 1988 13152
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12046
box 2340 12046 2540 12122
use cut_M2M3_1x2 
transform 1 0 1912 0 1 11984
box 1912 11984 1988 12184
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17242
box 2340 17242 2540 17318
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17180
box 1732 17180 1808 17380
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19662
box 2340 19662 2540 19738
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19600
box 1732 19600 1808 19800
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18210
box 2340 18210 2540 18286
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18148
box 1732 18148 1808 18348
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19178
box 2340 19178 2540 19254
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19116
box 1732 19116 1808 19316
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18694
box 2340 18694 2540 18770
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18632
box 1732 18632 1808 18832
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17726
box 2340 17726 2540 17802
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17664
box 1732 17664 1808 17864
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17242
box 2340 17242 2540 17318
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17180
box 1732 17180 1808 17380
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19662
box 2340 19662 2540 19738
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19600
box 1732 19600 1808 19800
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18210
box 2340 18210 2540 18286
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18148
box 1732 18148 1808 18348
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19178
box 2340 19178 2540 19254
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19116
box 1732 19116 1808 19316
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18694
box 2340 18694 2540 18770
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18632
box 1732 18632 1808 18832
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17726
box 2340 17726 2540 17802
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17664
box 1732 17664 1808 17864
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17242
box 2340 17242 2540 17318
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17180
box 1732 17180 1808 17380
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19662
box 2340 19662 2540 19738
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19600
box 1732 19600 1808 19800
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18210
box 2340 18210 2540 18286
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18148
box 1732 18148 1808 18348
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19178
box 2340 19178 2540 19254
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19116
box 1732 19116 1808 19316
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18694
box 2340 18694 2540 18770
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18632
box 1732 18632 1808 18832
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17726
box 2340 17726 2540 17802
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17664
box 1732 17664 1808 17864
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17242
box 2340 17242 2540 17318
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17180
box 1732 17180 1808 17380
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19662
box 2340 19662 2540 19738
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19600
box 1732 19600 1808 19800
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18210
box 2340 18210 2540 18286
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18148
box 1732 18148 1808 18348
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19178
box 2340 19178 2540 19254
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19116
box 1732 19116 1808 19316
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18694
box 2340 18694 2540 18770
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18632
box 1732 18632 1808 18832
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17726
box 2340 17726 2540 17802
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17664
box 1732 17664 1808 17864
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17242
box 2340 17242 2540 17318
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17180
box 1732 17180 1808 17380
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19662
box 2340 19662 2540 19738
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19600
box 1732 19600 1808 19800
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18210
box 2340 18210 2540 18286
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18148
box 1732 18148 1808 18348
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19178
box 2340 19178 2540 19254
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19116
box 1732 19116 1808 19316
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18694
box 2340 18694 2540 18770
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18632
box 1732 18632 1808 18832
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17726
box 2340 17726 2540 17802
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17664
box 1732 17664 1808 17864
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17242
box 2340 17242 2540 17318
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17180
box 1732 17180 1808 17380
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19662
box 2340 19662 2540 19738
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19600
box 1732 19600 1808 19800
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18210
box 2340 18210 2540 18286
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18148
box 1732 18148 1808 18348
use cut_M1M3_2x1 
transform 1 0 2340 0 1 19178
box 2340 19178 2540 19254
use cut_M2M3_1x2 
transform 1 0 1732 0 1 19116
box 1732 19116 1808 19316
use cut_M1M3_2x1 
transform 1 0 2340 0 1 18694
box 2340 18694 2540 18770
use cut_M2M3_1x2 
transform 1 0 1732 0 1 18632
box 1732 18632 1808 18832
use cut_M1M3_2x1 
transform 1 0 2340 0 1 17726
box 2340 17726 2540 17802
use cut_M2M3_1x2 
transform 1 0 1732 0 1 17664
box 1732 17664 1808 17864
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3042
box 2340 3042 2540 3118
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2980
box 1552 2980 1628 3180
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5462
box 2340 5462 2540 5538
use cut_M2M3_1x2 
transform 1 0 1552 0 1 5400
box 1552 5400 1628 5600
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4010
box 2340 4010 2540 4086
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3948
box 1552 3948 1628 4148
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4978
box 2340 4978 2540 5054
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4916
box 1552 4916 1628 5116
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4494
box 2340 4494 2540 4570
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4432
box 1552 4432 1628 4632
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3526
box 2340 3526 2540 3602
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3464
box 1552 3464 1628 3664
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3042
box 2340 3042 2540 3118
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2980
box 1552 2980 1628 3180
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5462
box 2340 5462 2540 5538
use cut_M2M3_1x2 
transform 1 0 1552 0 1 5400
box 1552 5400 1628 5600
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4010
box 2340 4010 2540 4086
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3948
box 1552 3948 1628 4148
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4978
box 2340 4978 2540 5054
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4916
box 1552 4916 1628 5116
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4494
box 2340 4494 2540 4570
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4432
box 1552 4432 1628 4632
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3526
box 2340 3526 2540 3602
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3464
box 1552 3464 1628 3664
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3042
box 2340 3042 2540 3118
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2980
box 1552 2980 1628 3180
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5462
box 2340 5462 2540 5538
use cut_M2M3_1x2 
transform 1 0 1552 0 1 5400
box 1552 5400 1628 5600
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4010
box 2340 4010 2540 4086
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3948
box 1552 3948 1628 4148
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4978
box 2340 4978 2540 5054
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4916
box 1552 4916 1628 5116
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4494
box 2340 4494 2540 4570
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4432
box 1552 4432 1628 4632
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3526
box 2340 3526 2540 3602
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3464
box 1552 3464 1628 3664
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3042
box 2340 3042 2540 3118
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2980
box 1552 2980 1628 3180
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5462
box 2340 5462 2540 5538
use cut_M2M3_1x2 
transform 1 0 1552 0 1 5400
box 1552 5400 1628 5600
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4010
box 2340 4010 2540 4086
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3948
box 1552 3948 1628 4148
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4978
box 2340 4978 2540 5054
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4916
box 1552 4916 1628 5116
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4494
box 2340 4494 2540 4570
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4432
box 1552 4432 1628 4632
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3526
box 2340 3526 2540 3602
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3464
box 1552 3464 1628 3664
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3042
box 2340 3042 2540 3118
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2980
box 1552 2980 1628 3180
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5462
box 2340 5462 2540 5538
use cut_M2M3_1x2 
transform 1 0 1552 0 1 5400
box 1552 5400 1628 5600
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4010
box 2340 4010 2540 4086
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3948
box 1552 3948 1628 4148
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4978
box 2340 4978 2540 5054
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4916
box 1552 4916 1628 5116
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4494
box 2340 4494 2540 4570
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4432
box 1552 4432 1628 4632
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3526
box 2340 3526 2540 3602
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3464
box 1552 3464 1628 3664
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3042
box 2340 3042 2540 3118
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2980
box 1552 2980 1628 3180
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5462
box 2340 5462 2540 5538
use cut_M2M3_1x2 
transform 1 0 1552 0 1 5400
box 1552 5400 1628 5600
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4010
box 2340 4010 2540 4086
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3948
box 1552 3948 1628 4148
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4978
box 2340 4978 2540 5054
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4916
box 1552 4916 1628 5116
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4494
box 2340 4494 2540 4570
use cut_M2M3_1x2 
transform 1 0 1552 0 1 4432
box 1552 4432 1628 4632
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3526
box 2340 3526 2540 3602
use cut_M2M3_1x2 
transform 1 0 1552 0 1 3464
box 1552 3464 1628 3664
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6366
box 2340 6366 2540 6442
use cut_M2M3_1x2 
transform 1 0 1372 0 1 6304
box 1372 6304 1448 6504
use cut_M1M3_2x1 
transform 1 0 2340 0 1 14886
box 2340 14886 2540 14962
use cut_M2M3_1x2 
transform 1 0 1192 0 1 14824
box 1192 14824 1268 15024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 14402
box 2340 14402 2540 14478
use cut_M2M3_1x2 
transform 1 0 1012 0 1 14340
box 1012 14340 1088 14540
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16822
box 2340 16822 2540 16898
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16760
box 1012 16760 1088 16960
use cut_M1M3_2x1 
transform 1 0 2340 0 1 15370
box 2340 15370 2540 15446
use cut_M2M3_1x2 
transform 1 0 1012 0 1 15308
box 1012 15308 1088 15508
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16338
box 2340 16338 2540 16414
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16276
box 1012 16276 1088 16476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 14402
box 2340 14402 2540 14478
use cut_M2M3_1x2 
transform 1 0 1012 0 1 14340
box 1012 14340 1088 14540
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16822
box 2340 16822 2540 16898
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16760
box 1012 16760 1088 16960
use cut_M1M3_2x1 
transform 1 0 2340 0 1 15370
box 2340 15370 2540 15446
use cut_M2M3_1x2 
transform 1 0 1012 0 1 15308
box 1012 15308 1088 15508
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16338
box 2340 16338 2540 16414
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16276
box 1012 16276 1088 16476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 14402
box 2340 14402 2540 14478
use cut_M2M3_1x2 
transform 1 0 1012 0 1 14340
box 1012 14340 1088 14540
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16822
box 2340 16822 2540 16898
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16760
box 1012 16760 1088 16960
use cut_M1M3_2x1 
transform 1 0 2340 0 1 15370
box 2340 15370 2540 15446
use cut_M2M3_1x2 
transform 1 0 1012 0 1 15308
box 1012 15308 1088 15508
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16338
box 2340 16338 2540 16414
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16276
box 1012 16276 1088 16476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 14402
box 2340 14402 2540 14478
use cut_M2M3_1x2 
transform 1 0 1012 0 1 14340
box 1012 14340 1088 14540
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16822
box 2340 16822 2540 16898
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16760
box 1012 16760 1088 16960
use cut_M1M3_2x1 
transform 1 0 2340 0 1 15370
box 2340 15370 2540 15446
use cut_M2M3_1x2 
transform 1 0 1012 0 1 15308
box 1012 15308 1088 15508
use cut_M1M3_2x1 
transform 1 0 2340 0 1 16338
box 2340 16338 2540 16414
use cut_M2M3_1x2 
transform 1 0 1012 0 1 16276
box 1012 16276 1088 16476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 15854
box 2340 15854 2540 15930
use cut_M2M3_1x2 
transform 1 0 832 0 1 15792
box 832 15792 908 15992
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7334
box 2340 7334 2540 7410
use cut_M2M3_1x2 
transform 1 0 652 0 1 7272
box 652 7272 728 7472
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7818
box 2340 7818 2540 7894
use cut_M2M3_1x2 
transform 1 0 472 0 1 7756
box 472 7756 548 7956
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6850
box 2340 6850 2540 6926
use cut_M2M3_1x2 
transform 1 0 292 0 1 6788
box 292 6788 368 6988
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8302
box 2340 8302 2540 8378
use cut_M2M3_1x2 
transform 1 0 112 0 1 8240
box 112 8240 188 8440
use cut_M1M2_1x2 
transform 1 0 2668 0 1 5828
box 2668 5828 2736 6012
use cut_M1M2_1x2 
transform 1 0 2668 0 1 5828
box 2668 5828 2736 6012
<< labels >>
flabel m1 s 2100 8660 2160 22720 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew
flabel m1 s 1920 140 1980 22720 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew
flabel m1 s 1740 17180 1800 22720 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew
flabel m1 s 1560 2980 1620 22720 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew
flabel m1 s 1380 6304 1440 22720 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew
flabel m1 s 1200 14824 1260 22720 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew
flabel m1 s 1020 14340 1080 22720 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew
flabel m1 s 840 15792 900 22720 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew
flabel m1 s 660 7272 720 22720 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew
flabel m1 s 480 7756 540 22720 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew
flabel m1 s 300 6788 360 22720 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew
flabel m1 s 120 8240 180 22720 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew
flabel m1 s 2668 0 11768 76 0 FreeSans 400 0 0 0 AVSS
port 14 nsew
flabel m3 s 2668 19880 2744 22780 0 FreeSans 400 0 0 0 CTOP
port 13 nsew
<< end >>
