magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 2028 18720
<< locali >>
rect 1788 0 2028 18720
rect 0 0 2028 240
rect 0 18480 2028 18720
rect 0 0 240 18720
rect 1788 0 2028 18720
rect 816 530 984 590
rect 984 530 1044 590
rect 1020 678 1200 738
rect 1020 2378 1248 2438
rect 816 882 1020 942
rect 1020 4138 1248 4198
rect 816 2642 1020 2702
rect 1020 5898 1248 5958
rect 816 4402 1020 4462
rect 1020 7658 1248 7718
rect 816 6162 1020 6222
rect 1020 9418 1248 9478
rect 816 7922 1020 7982
rect 1020 11178 1248 11238
rect 816 9682 1020 9742
rect 1020 12938 1248 12998
rect 816 11442 1020 11502
rect 1020 14698 1248 14758
rect 816 13202 1020 13262
rect 1020 16458 1248 16518
rect 816 14962 1020 15022
rect 1020 18218 1248 18278
rect 816 16722 1020 16782
rect 1020 678 1080 18278
rect 1140 618 1248 678
rect 1356 442 2028 502
rect 1356 794 2028 854
rect 1356 2554 2028 2614
rect 1356 4314 2028 4374
rect 1356 6074 2028 6134
rect 1356 7834 2028 7894
rect 1356 9594 2028 9654
rect 1356 11354 2028 11414
rect 1356 13114 2028 13174
rect 1356 14874 2028 14934
rect 1356 16634 2028 16694
rect 0 516 276 576
rect 0 868 276 928
rect 0 2628 276 2688
rect 0 4388 276 4448
rect 0 6148 276 6208
rect 0 7908 276 7968
rect 0 9668 276 9728
rect 0 11428 276 11488
rect 0 13188 276 13248
rect 0 14948 276 15008
rect 0 16708 276 16768
<< m2 >>
rect 1812 618 2028 678
rect 0 530 216 590
rect 1812 618 2028 678
rect 1000 618 1248 694
rect 1000 618 1920 694
rect 1000 618 1076 694
rect 0 530 216 590
rect 568 530 816 606
rect 108 530 568 606
rect 568 530 644 606
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa20
transform 1 0 384 0 1 384
box 384 384 1644 736
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa30
transform 1 0 384 0 1 736
box 384 736 1644 2496
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa31
transform 1 0 384 0 1 2496
box 384 2496 1644 4256
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa32
transform 1 0 384 0 1 4256
box 384 4256 1644 6016
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa33
transform 1 0 384 0 1 6016
box 384 6016 1644 7776
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa34
transform 1 0 384 0 1 7776
box 384 7776 1644 9536
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa35
transform 1 0 384 0 1 9536
box 384 9536 1644 11296
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa36
transform 1 0 384 0 1 11296
box 384 11296 1644 13056
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa37
transform 1 0 384 0 1 13056
box 384 13056 1644 14816
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa38
transform 1 0 384 0 1 14816
box 384 14816 1644 16576
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa39
transform 1 0 384 0 1 16576
box 384 16576 1644 18336
use cut_M1M3_2x1 
transform 1 0 1156 0 1 618
box 1156 618 1356 694
use cut_M1M3_2x1 
transform 1 0 724 0 1 530
box 724 530 924 606
<< labels >>
flabel locali s 1788 0 2028 18720 0 FreeSans 400 0 0 0 AVSS
port 3 nsew
flabel m2 s 1812 618 2028 678 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew
flabel m2 s 0 530 216 590 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 2 nsew
<< end >>
