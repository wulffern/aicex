magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 1280
<< locali >>
rect 1230 530 1290 750
rect 1230 850 1290 1070
rect 720 210 858 270
rect 720 530 858 590
rect 720 690 858 750
rect 858 210 918 750
rect 1062 370 1260 430
rect 720 1170 1062 1230
rect 1062 370 1122 1230
rect 1260 50 1398 110
rect 1398 1090 1620 1150
rect 1398 50 1458 1150
rect 630 50 1350 110
<< poly >>
rect 270 462 1710 498
rect 270 782 1710 818
rect 270 1102 1710 1138
<< m3 >>
rect 1170 0 1354 1280
rect 630 0 814 1280
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 990 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 990 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 990 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 990 1280
use PCHDL MP0
transform 1 0 990 0 1 0
box 990 0 1980 320
use PCHDL MP1
transform 1 0 990 0 1 320
box 990 320 1980 640
use PCHDL MP2
transform 1 0 990 0 1 640
box 990 640 1980 960
use PCHDL MP3
transform 1 0 990 0 1 960
box 990 960 1980 1280
use cut_M1M4_2x1 
transform 1 0 1170 0 1 210
box 1170 210 1354 278
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1170
box 1170 1170 1354 1238
use cut_M1M4_2x1 
transform 1 0 630 0 1 370
box 630 370 814 438
use cut_M1M4_2x1 
transform 1 0 630 0 1 850
box 630 850 814 918
use cut_M1M4_2x1 
transform 1 0 630 0 1 1010
box 630 1010 814 1078
<< labels >>
flabel locali s 1890 120 2070 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 270 770 450 830 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 1530 130 1710 190 0 FreeSans 400 0 0 0 RST_N
port 5 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 EN
port 6 nsew
flabel locali s 1170 370 1350 430 0 FreeSans 400 0 0 0 ENO
port 7 nsew
flabel m3 s 1170 0 1354 1280 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 1280 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
