magic
tech sky130A
magscale 1 2
timestamp 1661983200
<< checkpaint >>
rect 0 0 48580 63440
<< locali >>
rect 47812 528 48052 62912
rect 528 528 48052 768
rect 528 62672 48052 62912
rect 528 528 768 62912
rect 47812 528 48052 62912
rect 48340 0 48580 63440
rect 0 0 48580 240
rect 0 63200 48580 63440
rect 0 0 240 63440
rect 48340 0 48580 63440
rect 18568 8016 32704 8076
<< m2 >>
rect 41080 24754 41296 24814
rect 1056 1970 1272 2030
<< m1 >>
rect 29740 1056 29956 1116
use SUN_PLL_BUF xb1
transform 1 0 1056 0 1 1056
box 1056 1056 15768 12096
use SUN_PLL_LPF xb2
transform 1 0 1056 0 1 12536
box 1056 12536 40888 62384
use SUN_PLL_DIVN xc1
transform 1 0 18568 0 1 1056
box 18568 1056 32704 8092
use SUN_PLL_ROSC xd1
transform 1 0 33064 0 1 1056
box 33064 1056 39640 6464
use SUN_PLL_KICK xk1
transform 1 0 41080 0 1 1056
box 41080 1056 45208 11568
use SUN_PLL_CP xk2
transform 1 0 41080 0 1 12008
box 41080 12008 45496 22696
use SUN_PLL_PFD xk3
transform 1 0 41080 0 1 23136
box 41080 23136 45136 28896
use SUN_PLL_BIAS xl1
transform 1 0 45496 0 1 1056
box 45496 1056 47524 19776
<< labels >>
flabel locali s 47812 528 48052 62912 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 48340 0 48580 63440 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 18568 8016 32704 8076 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel m2 s 41080 24754 41296 24814 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel m1 s 29740 1056 29956 1116 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel m2 s 1056 1970 1272 2030 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
