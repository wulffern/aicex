magic
tech sky130A
magscale 1 2
timestamp 1659811303
<< checkpaint >>
rect 0 0 2520 704
<< locali >>
rect 432 498 600 558
rect 600 58 864 118
rect 600 58 660 558
rect 864 58 1032 118
rect 1032 58 1656 118
rect 1032 58 1092 118
rect 864 586 1032 646
rect 1032 586 1656 646
rect 1032 586 1092 646
rect 324 146 540 206
rect 756 586 972 646
<< poly >>
rect 324 158 2196 194
rect 324 510 2196 546
<< m3 >>
rect 1548 0 1748 704
rect 756 0 956 704
rect 1548 0 1748 704
rect 756 0 956 704
use SUNTR_NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_NCHDL MN1
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTR_PCHDL MP0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTR_PCHDL MP1
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTR_cut_M1M4_2x1 
transform 1 0 1548 0 1 234
box 1548 234 1748 310
use SUNTR_cut_M1M4_2x1 
transform 1 0 1548 0 1 410
box 1548 410 1748 486
use SUNTR_cut_M1M4_2x1 
transform 1 0 756 0 1 234
box 756 234 956 310
use SUNTR_cut_M1M4_2x1 
transform 1 0 756 0 1 410
box 756 410 956 486
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 756 586 972 646 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel m3 s 1548 0 1748 704 0 FreeSans 400 0 0 0 AVDD
port 3 nsew
flabel m3 s 756 0 956 704 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
<< end >>
