*RPLY_TEMP_SKY130A/RPLYTEMP_BG


*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLYTEMP_BG_lpe.spi
#else
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_10_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_20_lpe.spi
*.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_1_lpe.spi
.include ../../../work/xsch/RPLYTEMP_BG.spice
#endif



*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12
#else
.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VPWR  PWRUP_1V8  VSS  pwl 0 0 20n 0 20.1n {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS PWRUP_1V8 LPO LPO IBP_1U RPLYTEMP_BG

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

V1 IBP_1U 0 dc {AVDD/2}

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.measure tran ibp_1u FIND i(V1) AT=100n


#ifdef Debug
.save all
#else
.probe v(VDD_1V8) v(VSS) v(PWRUP_1V8) v(LPI) v(LPO) v(IBP_1U) i(v1) v(XDUT.VD1) v(XDUT.VD2)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

#ifdef Debug
tran 1n 200n 1n
write
*quit
#else
tran 1n 200n 1n
write
quit
#endif

.endc

.end


