magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 2560
<< locali >>
rect 720 210 858 270
rect 720 370 858 430
rect 720 850 858 910
rect 720 1010 858 1070
rect 720 1490 858 1550
rect 720 1650 858 1710
rect 720 2130 858 2190
rect 720 2290 858 2350
rect 858 210 1260 270
rect 858 370 1260 430
rect 858 850 1260 910
rect 858 1010 1260 1070
rect 858 1490 1260 1550
rect 858 1650 1260 1710
rect 858 2130 1260 2190
rect 858 2290 1260 2350
rect 858 210 918 2350
rect 330 130 390 2430
rect 1590 130 1650 2430
<< poly >>
rect 270 142 1710 178
rect 270 462 1710 498
rect 270 782 1710 818
rect 270 1102 1710 1138
rect 270 1422 1710 1458
rect 270 1742 1710 1778
rect 270 2062 1710 2098
rect 270 2382 1710 2418
<< m3 >>
rect 1170 0 1354 2560
rect 630 0 814 2560
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 990 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 990 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 990 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 990 1280
use NCHDL MN4
transform 1 0 0 0 1 1280
box 0 1280 990 1600
use NCHDL MN5
transform 1 0 0 0 1 1600
box 0 1600 990 1920
use NCHDL MN6
transform 1 0 0 0 1 1920
box 0 1920 990 2240
use NCHDL MN7
transform 1 0 0 0 1 2240
box 0 2240 990 2560
use PCHDL MP0
transform 1 0 990 0 1 0
box 990 0 1980 320
use PCHDL MP1
transform 1 0 990 0 1 320
box 990 320 1980 640
use PCHDL MP2
transform 1 0 990 0 1 640
box 990 640 1980 960
use PCHDL MP3
transform 1 0 990 0 1 960
box 990 960 1980 1280
use PCHDL MP4
transform 1 0 990 0 1 1280
box 990 1280 1980 1600
use PCHDL MP5
transform 1 0 990 0 1 1600
box 990 1600 1980 1920
use PCHDL MP6
transform 1 0 990 0 1 1920
box 990 1920 1980 2240
use PCHDL MP7
transform 1 0 990 0 1 2240
box 990 2240 1980 2560
use cut_M1M4_2x1 
transform 1 0 1170 0 1 50
box 1170 50 1354 118
use cut_M1M4_2x1 
transform 1 0 1170 0 1 530
box 1170 530 1354 598
use cut_M1M4_2x1 
transform 1 0 1170 0 1 690
box 1170 690 1354 758
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1170
box 1170 1170 1354 1238
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1330
box 1170 1330 1354 1398
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1810
box 1170 1810 1354 1878
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1970
box 1170 1970 1354 2038
use cut_M1M4_2x1 
transform 1 0 1170 0 1 2450
box 1170 2450 1354 2518
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M4_2x1 
transform 1 0 630 0 1 690
box 630 690 814 758
use cut_M1M4_2x1 
transform 1 0 630 0 1 1170
box 630 1170 814 1238
use cut_M1M4_2x1 
transform 1 0 630 0 1 1330
box 630 1330 814 1398
use cut_M1M4_2x1 
transform 1 0 630 0 1 1810
box 630 1810 814 1878
use cut_M1M4_2x1 
transform 1 0 630 0 1 1970
box 630 1970 814 2038
use cut_M1M4_2x1 
transform 1 0 630 0 1 2450
box 630 2450 814 2518
<< labels >>
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 630 210 810 270 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel locali s 1890 120 2070 200 0 FreeSans 400 0 0 0 BULKP
port 3 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 4 nsew
flabel m3 s 1170 0 1354 2560 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 630 0 814 2560 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
