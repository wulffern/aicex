magic
tech sky130A
magscale 1 2
timestamp 1660664629
<< checkpaint >>
rect 0 0 200 200
<< locali >>
rect 0 0 184 184
<< m1 >>
rect 0 0 184 184
<< m2 >>
rect 0 0 200 200
<< m3 >>
rect 0 0 200 200
<< viali >>
rect 12 12 172 172
<< v1 >>
rect 12 12 172 172
<< v2 >>
rect 12 12 188 188
<< labels >>
<< end >>
