**********************************************************************
**        Copyright (c) 2016 Carsten Wulff Software, Norway
** *******************************************************************
** Created       : wulff at 2016-11-16
** *******************************************************************

*-----------------------------------------------------------------------------
* Inverters
*-----------------------------------------------------------------------------

.subckt TIEH_CV Y  AVDD AVSS
MN0 A A AVSS AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
.ends

.subckt TIEL_CV Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 A A AVDD AVDD PCHDL
.ends TIEL_CV


.subckt IVX1_CV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
.ends

.subckt IVX2_CV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
MP1 AVDD A Y AVDD PCHDL
.ends

.subckt IVX4_CV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
MP1 AVDD A Y AVDD PCHDL
MP2 Y A AVDD AVDD PCHDL
MP3 AVDD A Y AVDD PCHDL
.ends IVX4_CV

.subckt IVX8_CV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MN4 Y A AVSS AVSS NCHDL
MN5 AVSS A Y AVSS NCHDL
MN6 Y A AVSS AVSS NCHDL
MN7 AVSS A Y AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
MP1 AVDD A Y AVDD PCHDL
MP2 Y A AVDD AVDD PCHDL
MP3 AVDD A Y AVDD PCHDL
MP4 Y A AVDD AVDD PCHDL
MP5 AVDD A Y AVDD PCHDL
MP6 Y A AVDD AVDD PCHDL
MP7 AVDD A Y AVDD PCHDL
.ends IVX8_CV

*-----------------------------------------------------------------------------
* Buffer
*-----------------------------------------------------------------------------

.subckt BFX1_CV A Y AVDD AVSS
MN0 AVSS A B AVSS NCHDL
MN1 Y B AVSS AVSS NCHDL
MP0 AVDD A B AVDD PCHDL
MP1 Y B AVDD AVDD PCHDL
.ends BFX1_CV



*-----------------------------------------------------------------------------
* NAND/NOR
*-----------------------------------------------------------------------------

.subckt NRX1_CV A B Y AVDD AVSS
MN0 Y A AVSS AVSS  NCHDL
MN1 AVSS B Y AVSS  NCHDL
MP0 N1 A AVDD AVDD PCHDL
MP1 Y B N1 AVDD PCHDL
.ends NRX1_CV

.subckt NDX1_CV A B Y AVDD AVSS
MN0 N1 A AVSS AVSS NCHDL
MN1 Y B N1 AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
MP1 AVDD B Y AVDD PCHDL
.ends NDX1_CV

.subckt ORX1_CV A B Y  AVDD AVSS
XA1 A B YN  AVDD AVSS  NRX1_CV
XA2 YN Y  AVDD AVSS  IVX1_CV
.ends

.subckt ANX1_CV A B Y  AVDD AVSS
XA1 A B YN  AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ends


.subckt IVTRIX1_CV A C CN Y AVDD AVSS
MN0 N1 A AVSS AVSS NCHDL
MN1 Y C N1 AVSS NCHDL
MP0 N2 A AVDD AVDD PCHDL
MP1 Y CN N2 AVDD PCHDL
.ends IVTRIX1_CV

.subckt NDTRIX1_CV A C CN RN Y AVDD AVSS
MN2 N1 RN AVSS AVSS NCHDL
MN0 N2 A N1 AVSS NCHDL
MN1 Y C N2 AVSS NCHDL
MP2 AVDD RN N2 AVDD PCHDL
MP0 N2 A AVDD AVDD PCHDL
MP1 Y CN N2 AVDD PCHDL
.ends

.subckt NRTRIX1_CV A C CN B Y AVDD AVSS
MN2 N1 B AVSS AVSS NCHDL
MN0 AVSS A N1 AVSS NCHDL
MN1 N1 C Y AVSS NCHDL
MP2 N2 B AVDD AVDD PCHDL
MP0 AVDD A N2 AVDD PCHDL
MP1 N2 CN Y AVDD PCHDL
.ends


.subckt DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS IVX1_CV
XA3 D CKN CKB A0  AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0  AVDD AVSS IVTRIX1_CV
XA5 A0 A1  AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN  AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN  AVDD AVSS NDTRIX1_CV
XA8 QN Q  AVDD AVSS IVX1_CV
.ends


.SUBCKT SCX1_CV A Y  AVDD AVSS
XA2 N1 A AVSS AVSS  NCHDL
XA3 SCO A N1 AVSS  NCHDL
XA4a AVDD SCO N1 AVSS  NCHDL
XA4b AVDD SCO N1 AVSS  NCHDL
XA5 Y SCO AVSS AVSS  NCHDL

XB0 N2 A AVDD AVDD  PCHDL
XB1 SCO A N2 AVDD  PCHDL
XB3a N2 SCO AVSS AVDD  PCHDL
XB3b N2 SCO AVSS AVDD  PCHDL
XB4 Y SCO AVDD AVDD  PCHDL
.ends




.SUBCKT TAPCELLB_CV AVDD AVSS
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 AVDD AVDD AVDD AVDD  PCHDL
.ENDS


.subckt SWX2_CV A Y VREF AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVDD PCHDL
MP1 VREF A Y AVDD PCHDL
.ends SWX2_CV


.subckt SWX4_CV A Y VREF  AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVDD PCHDL
MP1 VREF A Y AVDD PCHDL
MP2 Y A VREF AVDD PCHDL
MP3 VREF A Y AVDD PCHDL
.ends IVX4_CV

.subckt TGPD_CV C A B  AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN1 B C AVSS AVSS NCHDL
MN2 A CN B AVSS NCHDL
MP0 AVDD C CN AVDD PCHDL
MP1_DMY B AVDD AVDD AVDD PCHDL
MP2 A C B AVDD PCHDL
.ends

.subckt DFTSPCX1_CV D CK Q AVDD AVSS
MN0 N1 D AVSS AVSS NCHDL
MN2 N2 CK Q AVSS NCHDL
MN1 AVSS N1 N2 AVSS NCHDL
MP1 N3 D AVDD AVDD PCHDL
MP0 N1 CK N3 AVDD PCHDL
MP2 Q N1 AVDD AVDD PCHDL
.ends


.subckt SUN_TR AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 Y1 AVDD AVSS TIEH_CV
XA2 Y2 AVDD AVSS TIEL_CV
XB0 AVDD AVSS TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS IVX1_CV
XB4 A4 Y4 AVDD AVSS IVX2_CV
XB5 A5 Y5 AVDD AVSS IVX4_CV
XB6 A6 Y6 AVDD AVSS IVX8_CV
XC0 AVDD AVSS TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS BFX1_CV
XD0 AVDD AVSS TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS ANX1_CV
XE0 AVDD AVSS TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SCX1_CV
XF0 AVDD AVSS TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS TGPD_CV
XF18 A16 B16 Y16 AVDD AVSS DFTSPCX1_CV
.ends
