*RPLY_BIAS_SKY130A/RPLYBS_OTA
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLYBS_OTA_lpe.spi
#else
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_10_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_20_lpe.spi
.include ../../../work/xsch/RPLYBS_OTA.spice
#endif

.include ../balun.spi

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
*.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12
#else
*.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param vcm = 0.6
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc {vdda}
VPWR PWRUP_1V8 0 dc {vdda}

VI VI 0 dc 1m ac 1
VC VC 0 dc {vcm}

XB VI VC VIP VIN balun

IB 0 IBP_2U dc 2u

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VO VSS PWRUP_1V8 VIN VIP IBP_2U RPLYBS_OTA

*----------------------------------------------------------------
* WAVES
*----------------------------------------------------------------


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------
.measure dc vcm2 FIND par('(v(xdut.vin_ls) + v(xdut.vip_ls))/2') AT={0}
.measure dc vs FIND v(xdut.vs) AT={0}
.measure dc vbn1 FIND v(xdut.vbn1) AT={0}
.measure dc vbn2 FIND v(xdut.vbn1) AT={0}


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save all
.probe v(VDD_1V8) v(VO) v(VSS) v(PWRUP_1V8) v(VIN) v(VIP) v(gain_large_db)
+ v(gain_small_db)
+ v(VI)
+ v(xdut.vbn1)
+ v(xdut.vbn2)
+ v(xdut.vs)
+ v(xdut.vin_ls)
+ v(xdut.vip_ls)
#endif


*.dc VI -{vcm} {vcm} 1.1m

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*- Use a step that does not hit 0 to avoid infinite large signal gain
dc VI -0.5 0.5 1.1m

let asdb = 20*log10(abs(deriv(v(vo))/deriv(vi)))
let aldb = 20*log10(abs(v(vo)/v(vi)))
meas dc a_small_db_0  find asdb at=0
meas dc a_large_db_0  find aldb at=0
meas dc a_small_db_max  max asdb
meas dc a_large_db_max  max aldb
write
quit


.endc

.end
