magic
tech sky130A
magscale 1 2
timestamp 1660215182
<< checkpaint >>
rect -640 -640 4744 3500
<< locali >>
rect -640 -640 4744 -528
rect -640 -640 4744 -528
rect -640 -640 -528 3500
rect -640 3388 4744 3500
rect 4632 -640 4744 3500
rect -640 -640 4744 -528
rect 3834 2750 4158 2970
rect -54 2750 270 2970
<< ptapc >>
rect -628 -640 -548 -560
rect -548 -640 -468 -560
rect -468 -640 -388 -560
rect -388 -640 -308 -560
rect -308 -640 -228 -560
rect -228 -640 -148 -560
rect -148 -640 -68 -560
rect -68 -640 12 -560
rect 12 -640 92 -560
rect 92 -640 172 -560
rect 172 -640 252 -560
rect 252 -640 332 -560
rect 332 -640 412 -560
rect 412 -640 492 -560
rect 492 -640 572 -560
rect 572 -640 652 -560
rect 652 -640 732 -560
rect 732 -640 812 -560
rect 812 -640 892 -560
rect 892 -640 972 -560
rect 972 -640 1052 -560
rect 1052 -640 1132 -560
rect 1132 -640 1212 -560
rect 1212 -640 1292 -560
rect 1292 -640 1372 -560
rect 1372 -640 1452 -560
rect 1452 -640 1532 -560
rect 1532 -640 1612 -560
rect 1612 -640 1692 -560
rect 1692 -640 1772 -560
rect 1772 -640 1852 -560
rect 1852 -640 1932 -560
rect 1932 -640 2012 -560
rect 2012 -640 2092 -560
rect 2092 -640 2172 -560
rect 2172 -640 2252 -560
rect 2252 -640 2332 -560
rect 2332 -640 2412 -560
rect 2412 -640 2492 -560
rect 2492 -640 2572 -560
rect 2572 -640 2652 -560
rect 2652 -640 2732 -560
rect 2732 -640 2812 -560
rect 2812 -640 2892 -560
rect 2892 -640 2972 -560
rect 2972 -640 3052 -560
rect 3052 -640 3132 -560
rect 3132 -640 3212 -560
rect 3212 -640 3292 -560
rect 3292 -640 3372 -560
rect 3372 -640 3452 -560
rect 3452 -640 3532 -560
rect 3532 -640 3612 -560
rect 3612 -640 3692 -560
rect 3692 -640 3772 -560
rect 3772 -640 3852 -560
rect 3852 -640 3932 -560
rect 3932 -640 4012 -560
rect 4012 -640 4092 -560
rect 4092 -640 4172 -560
rect 4172 -640 4252 -560
rect 4252 -640 4332 -560
rect 4332 -640 4412 -560
rect 4412 -640 4492 -560
rect 4492 -640 4572 -560
rect 4572 -640 4652 -560
rect 4652 -640 4732 -560
rect -640 -610 -560 -530
rect -640 -530 -560 -450
rect -640 -450 -560 -370
rect -640 -370 -560 -290
rect -640 -290 -560 -210
rect -640 -210 -560 -130
rect -640 -130 -560 -50
rect -640 -50 -560 30
rect -640 30 -560 110
rect -640 110 -560 190
rect -640 190 -560 270
rect -640 270 -560 350
rect -640 350 -560 430
rect -640 430 -560 510
rect -640 510 -560 590
rect -640 590 -560 670
rect -640 670 -560 750
rect -640 750 -560 830
rect -640 830 -560 910
rect -640 910 -560 990
rect -640 990 -560 1070
rect -640 1070 -560 1150
rect -640 1150 -560 1230
rect -640 1230 -560 1310
rect -640 1310 -560 1390
rect -640 1390 -560 1470
rect -640 1470 -560 1550
rect -640 1550 -560 1630
rect -640 1630 -560 1710
rect -640 1710 -560 1790
rect -640 1790 -560 1870
rect -640 1870 -560 1950
rect -640 1950 -560 2030
rect -640 2030 -560 2110
rect -640 2110 -560 2190
rect -640 2190 -560 2270
rect -640 2270 -560 2350
rect -640 2350 -560 2430
rect -640 2430 -560 2510
rect -640 2510 -560 2590
rect -640 2590 -560 2670
rect -640 2670 -560 2750
rect -640 2750 -560 2830
rect -640 2830 -560 2910
rect -640 2910 -560 2990
rect -640 2990 -560 3070
rect -640 3070 -560 3150
rect -640 3150 -560 3230
rect -640 3230 -560 3310
rect -640 3310 -560 3390
rect -640 3390 -560 3470
rect -628 3388 -548 3468
rect -548 3388 -468 3468
rect -468 3388 -388 3468
rect -388 3388 -308 3468
rect -308 3388 -228 3468
rect -228 3388 -148 3468
rect -148 3388 -68 3468
rect -68 3388 12 3468
rect 12 3388 92 3468
rect 92 3388 172 3468
rect 172 3388 252 3468
rect 252 3388 332 3468
rect 332 3388 412 3468
rect 412 3388 492 3468
rect 492 3388 572 3468
rect 572 3388 652 3468
rect 652 3388 732 3468
rect 732 3388 812 3468
rect 812 3388 892 3468
rect 892 3388 972 3468
rect 972 3388 1052 3468
rect 1052 3388 1132 3468
rect 1132 3388 1212 3468
rect 1212 3388 1292 3468
rect 1292 3388 1372 3468
rect 1372 3388 1452 3468
rect 1452 3388 1532 3468
rect 1532 3388 1612 3468
rect 1612 3388 1692 3468
rect 1692 3388 1772 3468
rect 1772 3388 1852 3468
rect 1852 3388 1932 3468
rect 1932 3388 2012 3468
rect 2012 3388 2092 3468
rect 2092 3388 2172 3468
rect 2172 3388 2252 3468
rect 2252 3388 2332 3468
rect 2332 3388 2412 3468
rect 2412 3388 2492 3468
rect 2492 3388 2572 3468
rect 2572 3388 2652 3468
rect 2652 3388 2732 3468
rect 2732 3388 2812 3468
rect 2812 3388 2892 3468
rect 2892 3388 2972 3468
rect 2972 3388 3052 3468
rect 3052 3388 3132 3468
rect 3132 3388 3212 3468
rect 3212 3388 3292 3468
rect 3292 3388 3372 3468
rect 3372 3388 3452 3468
rect 3452 3388 3532 3468
rect 3532 3388 3612 3468
rect 3612 3388 3692 3468
rect 3692 3388 3772 3468
rect 3772 3388 3852 3468
rect 3852 3388 3932 3468
rect 3932 3388 4012 3468
rect 4012 3388 4092 3468
rect 4092 3388 4172 3468
rect 4172 3388 4252 3468
rect 4252 3388 4332 3468
rect 4332 3388 4412 3468
rect 4412 3388 4492 3468
rect 4492 3388 4572 3468
rect 4572 3388 4652 3468
rect 4652 3388 4732 3468
rect 4632 -610 4712 -530
rect 4632 -530 4712 -450
rect 4632 -450 4712 -370
rect 4632 -370 4712 -290
rect 4632 -290 4712 -210
rect 4632 -210 4712 -130
rect 4632 -130 4712 -50
rect 4632 -50 4712 30
rect 4632 30 4712 110
rect 4632 110 4712 190
rect 4632 190 4712 270
rect 4632 270 4712 350
rect 4632 350 4712 430
rect 4632 430 4712 510
rect 4632 510 4712 590
rect 4632 590 4712 670
rect 4632 670 4712 750
rect 4632 750 4712 830
rect 4632 830 4712 910
rect 4632 910 4712 990
rect 4632 990 4712 1070
rect 4632 1070 4712 1150
rect 4632 1150 4712 1230
rect 4632 1230 4712 1310
rect 4632 1310 4712 1390
rect 4632 1390 4712 1470
rect 4632 1470 4712 1550
rect 4632 1550 4712 1630
rect 4632 1630 4712 1710
rect 4632 1710 4712 1790
rect 4632 1790 4712 1870
rect 4632 1870 4712 1950
rect 4632 1950 4712 2030
rect 4632 2030 4712 2110
rect 4632 2110 4712 2190
rect 4632 2190 4712 2270
rect 4632 2270 4712 2350
rect 4632 2350 4712 2430
rect 4632 2430 4712 2510
rect 4632 2510 4712 2590
rect 4632 2590 4712 2670
rect 4632 2670 4712 2750
rect 4632 2750 4712 2830
rect 4632 2830 4712 2910
rect 4632 2910 4712 2990
rect 4632 2990 4712 3070
rect 4632 3070 4712 3150
rect 4632 3150 4712 3230
rect 4632 3230 4712 3310
rect 4632 3310 4712 3390
rect 4632 3390 4712 3470
<< ptap >>
rect -640 -640 4744 -528
rect -640 -640 -528 3500
rect -640 3388 4744 3500
rect 4632 -640 4744 3500
use SUNTR_RES200 XA1
transform 1 0 0 0 1 0
box 0 0 4104 2860
<< labels >>
flabel locali s -640 -640 4744 -528 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 3834 2750 4158 2970 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s -54 2750 270 2970 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
