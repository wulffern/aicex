**********************************************************************
**        Copyright (c) 2016 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2016-11-16
** *******************************************************************


.subckt TIEH_CV Y BULKP BULKN AVDD AVSS
MN0 A A AVSS BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
.ends

.subckt TIEL_CV Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MP0 A A AVDD BULKP PCHDL
.ends TIEL_CV


.subckt IVX1_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
.ends

.subckt TIVX1_CV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 Y A AVDD AVDD PCHDL
.ends

.subckt IVX2_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
.ends

.subckt IVX4_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
MP2 Y A AVDD BULKP PCHDL
MP3 AVDD A Y BULKP PCHDL
.ends IVX4_CV

.subckt IVX8_CV A Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MN4 Y A AVSS BULKN NCHDL
MN5 AVSS A Y BULKN NCHDL
MN6 Y A AVSS BULKN NCHDL
MN7 AVSS A Y BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD A Y BULKP PCHDL
MP2 Y A AVDD BULKP PCHDL
MP3 AVDD A Y BULKP PCHDL
MP4 Y A AVDD BULKP PCHDL
MP5 AVDD A Y BULKP PCHDL
MP6 Y A AVDD BULKP PCHDL
MP7 AVDD A Y BULKP PCHDL
.ends IVX8_CV

.subckt BFX1_CV A Y BULKP BULKN AVDD AVSS
MN0 AVSS A B BULKN NCHDL
MN1 Y B AVSS BULKN NCHDL
MP0 AVDD A B BULKP PCHDL
MP1 Y B AVDD BULKP PCHDL
.ends BFX1_CV


*-----------------------------------------------------------------------------
* NAND/NOR
*-----------------------------------------------------------------------------

.subckt NRX1_CV A B Y BULKP BULKN AVDD AVSS
MN0 Y A AVSS BULKN  NCHDL
MN1 AVSS B Y BULKN  NCHDL
MP0 N1 A AVDD BULKP PCHDL
MP1 Y B N1 BULKP PCHDL
.ends NRX1_CV

.subckt NDX1_CV A B Y BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y B N1 BULKN NCHDL
MP0 Y A AVDD BULKP PCHDL
MP1 AVDD B Y BULKP PCHDL
.ends NDX1_CV

.subckt ORX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS  NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS  IVX1_CV
.ends

.subckt ANX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS IVX1_CV
.ends


.subckt IVTRIX1_CV A C CN Y  BULKP BULKN AVDD AVSS
MN0 N1 A AVSS BULKN NCHDL
MN1 Y C N1 BULKN NCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends IVTRIX1_CV

.subckt NDTRIX1_CV A C CN RN Y BULKP BULKN AVDD AVSS
MN2 N1 RN AVSS BULKN NCHDL
MN0 N2 A N1 BULKN NCHDL
MN1 Y C N2 BULKN NCHDL
MP2 AVDD RN N2 BULKP PCHDL
MP0 N2 A AVDD BULKP PCHDL
MP1 Y CN N2 BULKP PCHDL
.ends


.subckt DFRNQNX1_CV D CK RN Q QN BULKP BULKN AVDD AVSS
XA0 BULKP BULKN TAPCELLB_CV
XA1 CK RN CKN BULKP BULKN AVDD AVSS NDX1_CV
XA2 CKN CKB BULKP BULKN AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 BULKP BULKN AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 BULKP BULKN AVDD AVSS IVTRIX1_CV
XA5 A0 A1 BULKP BULKN AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN BULKP BULKN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN BULKP BULKN AVDD AVSS NDTRIX1_CV
XA8 QN Q BULKP BULKN AVDD AVSS IVX1_CV
.ends


.SUBCKT SCX1_CV A Y BULKP BULKN  AVDD AVSS
XA2 N1 A AVSS BULKN  NCHDL
XA3 SCO A N1 BULKN  NCHDL
XA4a AVDD SCO N1 BULKN  NCHDL
XA4b AVDD SCO N1 BULKN  NCHDL
XA5 Y SCO AVSS BULKN  NCHDL

XB0 N2 A AVDD BULKP  PCHDL
XB1 SCO A N2 BULKP  PCHDL
XB3a N2 SCO AVSS BULKP  PCHDL
XB3b N2 SCO AVSS BULKP  PCHDL
XB4 Y SCO AVDD AVSS  PCHDL
.ends


*-----------------------------------------------------------------------------
* SAR unit logic cells
*---------------------------------------------------------------------------


.SUBCKT TAPCELLB_CV AVDD AVSS
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 AVDD AVDD AVDD AVDD  PCHDL
.ENDS

.SUBCKT TAPCELLBAVSS_CV AVDD AVSS
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 NC1 NC1 NC1 AVDD  PCHDL
.ENDS


.subckt SWX2_CV A Y VREF AVSS BULKP BULKN
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MP0 Y A VREF BULKP PCHDL
MP1 VREF A Y BULKP PCHDL
.ends SWX2_CV


.subckt SWX4_CV A Y VREF AVSS BULKP BULKN
MN0 Y A AVSS BULKN NCHDL
MN1 AVSS A Y BULKN NCHDL
MN2 Y A AVSS BULKN NCHDL
MN3 AVSS A Y BULKN NCHDL
MP0 Y A VREF BULKP PCHDL
MP1 VREF A Y BULKP PCHDL
MP2 Y A VREF BULKP PCHDL
MP3 VREF A Y BULKP PCHDL
.ends IVX4_CV

.subckt TGPD_CV C A B BULKP BULKN AVDD AVSS
MN0 AVSS C CN BULKN NCHDL
MN1 B C AVSS BULKN NCHDL
MN2 A CN B BULKN NCHDL
MP0 AVDD C CN BULKP PCHDL
MP1_DMY B AVDD AVDD BULKP PCHDL
MP2 A C B BULKP PCHDL
.ends

