magic
tech sky130A
magscale 1 2
timestamp 1664582400
<< checkpaint >>
rect 0 0 2520 1760
<< locali >>
rect 864 234 1032 294
rect 864 410 1032 470
rect 864 762 1032 822
rect 864 1114 1032 1174
rect 1032 234 1092 1174
rect 1428 234 1656 294
rect 1428 410 1656 470
rect 1428 938 1656 998
rect 1428 1290 1656 1350
rect 1428 234 1488 1350
rect 402 146 462 558
rect 2088 850 2256 910
rect 1656 586 2256 646
rect 2088 1202 2256 1262
rect 2088 1554 2256 1614
rect 2256 586 2316 1614
rect 204 850 432 910
rect 204 586 864 646
rect 204 1202 432 1262
rect 204 1554 432 1614
rect 204 586 264 1614
rect 636 938 864 998
rect 636 1290 864 1350
rect 636 938 696 1350
rect 864 1642 1032 1702
rect 1032 1642 1656 1702
rect 1032 1642 1092 1702
rect 864 1290 1032 1350
rect 1032 1466 1656 1526
rect 1032 1290 1092 1526
rect 1656 762 1824 822
rect 1656 1114 1824 1174
rect 1824 762 1884 1174
rect 324 146 540 206
rect 756 1642 972 1702
<< m1 >>
rect 864 1466 1032 1526
rect 1032 1114 1656 1174
rect 1032 1114 1092 1526
rect 864 586 1032 646
rect 1032 586 1656 646
rect 1032 586 1092 646
<< poly >>
rect 324 158 2196 194
rect 324 510 2196 546
<< m3 >>
rect 1548 0 1748 1760
rect 756 0 956 1760
rect 1548 0 1748 1760
rect 756 0 956 1760
use SUNTRB_NCHDL XA2
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTRB_NCHDL XA3
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTRB_NCHDL XA4a
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNTRB_NCHDL XA4b
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNTRB_NCHDL XA5
transform 1 0 0 0 1 1408
box 0 1408 1260 1760
use SUNTRB_PCHDL XB0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTRB_PCHDL XB1
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTRB_PCHDL XB3a
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNTRB_PCHDL XB3b
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNTRB_PCHDL XB4
transform 1 0 1260 0 1 1408
box 1260 1408 2520 1760
use SUNTRB_cut_M1M2_2x1 
transform 1 0 756 0 1 1466
box 756 1466 940 1534
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1548 0 1 1114
box 1548 1114 1732 1182
use SUNTRB_cut_M1M2_2x1 
transform 1 0 756 0 1 586
box 756 586 940 654
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1548 0 1 586
box 1548 586 1732 654
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use SUNTRB_cut_M1M4_2x1 
transform 1 0 1548 0 1 1466
box 1548 1466 1748 1542
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 58
box 756 58 956 134
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 1466
box 756 1466 956 1542
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 756 1642 972 1702 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel m3 s 1548 0 1748 1760 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 756 0 956 1760 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
