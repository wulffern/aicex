magic
tech sky130A
magscale 1 2
timestamp 1658582973
<< checkpaint >>
rect 0 0 1512 1056
<< m1 >>
rect 108 -44 1476 44
rect 1404 44 1476 132
rect 108 132 1332 220
rect 1404 132 1476 220
rect 108 220 180 308
rect 1404 220 1476 308
rect 108 308 180 396
rect 252 308 1476 396
rect 108 396 180 484
rect 1404 396 1476 484
rect 108 484 1332 572
rect 1404 484 1476 572
rect 108 572 180 660
rect 1404 572 1476 660
rect 108 660 180 748
rect 252 660 1476 748
rect 108 748 180 836
rect 108 836 1476 924
<< m2 >>
rect 108 -44 1476 44
rect 1404 44 1476 132
rect 108 132 1332 220
rect 1404 132 1476 220
rect 108 220 180 308
rect 1404 220 1476 308
rect 108 308 180 396
rect 252 308 1476 396
rect 108 396 180 484
rect 1404 396 1476 484
rect 108 484 1332 572
rect 1404 484 1476 572
rect 108 572 180 660
rect 1404 572 1476 660
rect 108 660 180 748
rect 252 660 1476 748
rect 108 748 180 836
rect 108 836 1476 924
<< locali >>
rect 108 -44 1476 44
rect 1404 44 1476 132
rect 108 132 1332 220
rect 1404 132 1476 220
rect 108 220 180 308
rect 1404 220 1476 308
rect 108 308 180 396
rect 252 308 1476 396
rect 108 396 180 484
rect 1404 396 1476 484
rect 108 484 1332 572
rect 1404 484 1476 572
rect 108 572 180 660
rect 1404 572 1476 660
rect 108 660 180 748
rect 252 660 1476 748
rect 108 748 180 836
rect 108 836 1476 924
<< v1 >>
rect 1116 -35 1188 -26
rect 1116 -26 1188 -17
rect 1116 -17 1188 -8
rect 1116 -8 1188 0
rect 1116 0 1188 8
rect 1116 8 1188 17
rect 1116 17 1188 26
rect 1116 26 1188 35
rect 1188 -35 1260 -26
rect 1188 -26 1260 -17
rect 1188 -17 1260 -8
rect 1188 -8 1260 0
rect 1188 0 1260 8
rect 1188 8 1260 17
rect 1188 17 1260 26
rect 1188 26 1260 35
rect 1260 -35 1332 -26
rect 1260 -26 1332 -17
rect 1260 -17 1332 -8
rect 1260 -8 1332 0
rect 1260 0 1332 8
rect 1260 8 1332 17
rect 1260 17 1332 26
rect 1260 26 1332 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 1116 316 1188 325
rect 1116 325 1188 334
rect 1116 334 1188 343
rect 1116 343 1188 352
rect 1116 352 1188 360
rect 1116 360 1188 369
rect 1116 369 1188 378
rect 1116 378 1188 387
rect 1188 316 1260 325
rect 1188 325 1260 334
rect 1188 334 1260 343
rect 1188 343 1260 352
rect 1188 352 1260 360
rect 1188 360 1260 369
rect 1188 369 1260 378
rect 1188 378 1260 387
rect 1260 316 1332 325
rect 1260 325 1332 334
rect 1260 334 1332 343
rect 1260 343 1332 352
rect 1260 352 1332 360
rect 1260 360 1332 369
rect 1260 369 1332 378
rect 1260 378 1332 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 1116 668 1188 677
rect 1116 677 1188 686
rect 1116 686 1188 695
rect 1116 695 1188 704
rect 1116 704 1188 712
rect 1116 712 1188 721
rect 1116 721 1188 730
rect 1116 730 1188 739
rect 1188 668 1260 677
rect 1188 677 1260 686
rect 1188 686 1260 695
rect 1188 695 1260 704
rect 1188 704 1260 712
rect 1188 712 1260 721
rect 1188 721 1260 730
rect 1188 730 1260 739
rect 1260 668 1332 677
rect 1260 677 1332 686
rect 1260 686 1332 695
rect 1260 695 1332 704
rect 1260 704 1332 712
rect 1260 712 1332 721
rect 1260 721 1332 730
rect 1260 730 1332 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 1116 -35 1188 -26
rect 1116 -26 1188 -17
rect 1116 -17 1188 -8
rect 1116 -8 1188 0
rect 1116 0 1188 8
rect 1116 8 1188 17
rect 1116 17 1188 26
rect 1116 26 1188 35
rect 1188 -35 1260 -26
rect 1188 -26 1260 -17
rect 1188 -17 1260 -8
rect 1188 -8 1260 0
rect 1188 0 1260 8
rect 1188 8 1260 17
rect 1188 17 1260 26
rect 1188 26 1260 35
rect 1260 -35 1332 -26
rect 1260 -26 1332 -17
rect 1260 -17 1332 -8
rect 1260 -8 1332 0
rect 1260 0 1332 8
rect 1260 8 1332 17
rect 1260 17 1332 26
rect 1260 26 1332 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 1116 316 1188 325
rect 1116 325 1188 334
rect 1116 334 1188 343
rect 1116 343 1188 352
rect 1116 352 1188 360
rect 1116 360 1188 369
rect 1116 369 1188 378
rect 1116 378 1188 387
rect 1188 316 1260 325
rect 1188 325 1260 334
rect 1188 334 1260 343
rect 1188 343 1260 352
rect 1188 352 1260 360
rect 1188 360 1260 369
rect 1188 369 1260 378
rect 1188 378 1260 387
rect 1260 316 1332 325
rect 1260 325 1332 334
rect 1260 334 1332 343
rect 1260 343 1332 352
rect 1260 352 1332 360
rect 1260 360 1332 369
rect 1260 369 1332 378
rect 1260 378 1332 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 1116 668 1188 677
rect 1116 677 1188 686
rect 1116 686 1188 695
rect 1116 695 1188 704
rect 1116 704 1188 712
rect 1116 712 1188 721
rect 1116 721 1188 730
rect 1116 730 1188 739
rect 1188 668 1260 677
rect 1188 677 1260 686
rect 1188 686 1260 695
rect 1188 695 1260 704
rect 1188 704 1260 712
rect 1188 712 1260 721
rect 1188 721 1260 730
rect 1188 730 1260 739
rect 1260 668 1332 677
rect 1260 677 1332 686
rect 1260 686 1332 695
rect 1260 695 1332 704
rect 1260 704 1332 712
rect 1260 712 1332 721
rect 1260 721 1332 730
rect 1260 730 1332 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 1116 -35 1188 -26
rect 1116 -26 1188 -17
rect 1116 -17 1188 -8
rect 1116 -8 1188 0
rect 1116 0 1188 8
rect 1116 8 1188 17
rect 1116 17 1188 26
rect 1116 26 1188 35
rect 1188 -35 1260 -26
rect 1188 -26 1260 -17
rect 1188 -17 1260 -8
rect 1188 -8 1260 0
rect 1188 0 1260 8
rect 1188 8 1260 17
rect 1188 17 1260 26
rect 1188 26 1260 35
rect 1260 -35 1332 -26
rect 1260 -26 1332 -17
rect 1260 -17 1332 -8
rect 1260 -8 1332 0
rect 1260 0 1332 8
rect 1260 8 1332 17
rect 1260 17 1332 26
rect 1260 26 1332 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 1116 316 1188 325
rect 1116 325 1188 334
rect 1116 334 1188 343
rect 1116 343 1188 352
rect 1116 352 1188 360
rect 1116 360 1188 369
rect 1116 369 1188 378
rect 1116 378 1188 387
rect 1188 316 1260 325
rect 1188 325 1260 334
rect 1188 334 1260 343
rect 1188 343 1260 352
rect 1188 352 1260 360
rect 1188 360 1260 369
rect 1188 369 1260 378
rect 1188 378 1260 387
rect 1260 316 1332 325
rect 1260 325 1332 334
rect 1260 334 1332 343
rect 1260 343 1332 352
rect 1260 352 1332 360
rect 1260 360 1332 369
rect 1260 369 1332 378
rect 1260 378 1332 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 1116 668 1188 677
rect 1116 677 1188 686
rect 1116 686 1188 695
rect 1116 695 1188 704
rect 1116 704 1188 712
rect 1116 712 1188 721
rect 1116 721 1188 730
rect 1116 730 1188 739
rect 1188 668 1260 677
rect 1188 677 1260 686
rect 1188 686 1260 695
rect 1188 695 1260 704
rect 1188 704 1260 712
rect 1188 712 1260 721
rect 1188 721 1260 730
rect 1188 730 1260 739
rect 1260 668 1332 677
rect 1260 677 1332 686
rect 1260 686 1332 695
rect 1260 695 1332 704
rect 1260 704 1332 712
rect 1260 712 1332 721
rect 1260 721 1332 730
rect 1260 730 1332 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 1476 44
rect 108 -44 1476 44
rect 1404 44 1476 132
rect 108 132 1116 220
rect 1188 132 1332 220
rect 1404 132 1476 220
rect 108 220 180 308
rect 1404 220 1476 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 1476 396
rect 108 396 180 484
rect 1404 396 1476 484
rect 108 484 1332 572
rect 1404 484 1476 572
rect 108 572 180 660
rect 1404 572 1476 660
rect 108 660 180 748
rect 252 660 1476 748
rect 108 748 180 836
rect 108 836 1476 924
rect 108 836 1476 924
<< rm3 >>
rect 1116 132 1188 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 1476 44 0 FreeSans 400 0 0 0 B
port 1 nsew
flabel m3 s 108 836 1476 924 0 FreeSans 400 0 0 0 A
port 2 nsew
<< end >>
