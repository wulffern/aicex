
*-------------------------------------------------------------
* SUNPLL_SUNTR_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_NCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_NCHDLCM D G S B
XM0 N0 G S B SUNPLL_SUNTR_NCHDL
XM1 N1 G N0 B SUNPLL_SUNTR_NCHDL
XM2 N2 G N1 B SUNPLL_SUNTR_NCHDL
XM3 N3 G N2 B SUNPLL_SUNTR_NCHDL
XM4 N4 G N3 B SUNPLL_SUNTR_NCHDL
XM5 N5 G N4 B SUNPLL_SUNTR_NCHDL
XM6 N6 G N5 B SUNPLL_SUNTR_NCHDL
XM7 N7 G N6 B SUNPLL_SUNTR_NCHDL
XM8 D G N7 B SUNPLL_SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_PCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_PCHDLCM D G S B
XM0 N0 G S B SUNPLL_SUNTR_PCHDL
XM7 D G N0 B SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_NCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_NCHDLA D G S B
XM0 D G S B SUNPLL_SUNTR_NCHDL
XM1 S G D B SUNPLL_SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_PCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_PCHDLA D G S B
XM0 D G S B SUNPLL_SUNTR_PCHDL
XM1 S G D B SUNPLL_SUNTR_PCHDL
XM2 D G S B SUNPLL_SUNTR_PCHDL
XM3 S G D B SUNPLL_SUNTR_PCHDL
XM4 D G S B SUNPLL_SUNTR_PCHDL
XM5 S G D B SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_RES12 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_RES12 N P B
XRR1_0 N INT_0 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_1 INT_0 P B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_RPPO_12k <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_RPPO_12k P N B
XA1 N P B SUNPLL_SUNTR_RES12
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_TAPCELLB_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNPLL_SUNTR_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_IVX1_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNPLL_SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_NRX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_NRX1_CV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNPLL_SUNTR_NCHDL
XMN1 AVSS B Y AVSS SUNPLL_SUNTR_NCHDL
XMP0 N1 A AVDD AVDD SUNPLL_SUNTR_PCHDL
XMP1 Y B N1 AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_NDX1_CV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNPLL_SUNTR_NCHDL
XMN1 Y B N1 AVSS SUNPLL_SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNPLL_SUNTR_PCHDL
XMP1 AVDD B Y AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_DFTSPCX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_DFTSPCX1_CV D CK Q AVDD AVSS
XMN0 N1 D AVSS AVSS SUNPLL_SUNTR_NCHDL
XMN2 N2 CK Q AVSS SUNPLL_SUNTR_NCHDL
XMN1 AVSS N1 N2 AVSS SUNPLL_SUNTR_NCHDL
XMP1 N3 D AVDD AVDD SUNPLL_SUNTR_PCHDL
XMP0 N1 CK N3 AVDD SUNPLL_SUNTR_PCHDL
XMP2 Q N1 AVDD AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_IVTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_IVTRIX1_CV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNPLL_SUNTR_NCHDL
XMN1 Y C N1 AVSS SUNPLL_SUNTR_NCHDL
XMP0 N2 A AVDD AVDD SUNPLL_SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_NDTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_NDTRIX1_CV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS SUNPLL_SUNTR_NCHDL
XMN0 N2 A N1 AVSS SUNPLL_SUNTR_NCHDL
XMN1 Y C N2 AVSS SUNPLL_SUNTR_NCHDL
XMP2 AVDD RN N2 AVDD SUNPLL_SUNTR_PCHDL
XMP0 N2 A AVDD AVDD SUNPLL_SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTR_DFRNQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS SUNPLL_SUNTR_TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS SUNPLL_SUNTR_NDX1_CV
XA2 CKN CKB AVDD AVSS SUNPLL_SUNTR_IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS SUNPLL_SUNTR_IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS SUNPLL_SUNTR_IVTRIX1_CV
XA5 A0 A1 AVDD AVSS SUNPLL_SUNTR_IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS SUNPLL_SUNTR_IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS SUNPLL_SUNTR_NDTRIX1_CV
XA8 QN Q AVDD AVSS SUNPLL_SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTRB_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTRB_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTRB_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTRB_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTRB_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTRB_IVX1_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNPLL_SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNPLL_SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTRB_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTRB_NDX1_CV A B Y BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNPLL_SUNTRB_NCHDL
XMN1 Y B N1 BULKN SUNPLL_SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNPLL_SUNTRB_PCHDL
XMP1 AVDD B Y BULKP SUNPLL_SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNTRB_TAPCELLBAVSS_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNTRB_TAPCELLBAVSS_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNPLL_SUNTRB_NCHDL
XMP1 NC1 NC1 NC1 AVDD SUNPLL_SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUNSAR_CAP_BSSW_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUNSAR_CAP_BSSW_CV A B
RR1 A NC0 sky130_fd_pr__res_generic_m1  l=0.36  w=0.44  
RR2 B NC1 sky130_fd_pr__res_generic_m1  l=0.36  w=0.44  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_LSCORE <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_LSCORE A AN YN Y AVDD AVSS
xb1_0 Y AN AVSS AVSS SUNPLL_SUNTR_NCHDL
xb1_1 Y AN AVSS AVSS SUNPLL_SUNTR_NCHDL
xb2_0 YN A AVSS AVSS SUNPLL_SUNTR_NCHDL
xb2_1 YN A AVSS AVSS SUNPLL_SUNTR_NCHDL
xc1a net2 YN AVDD AVDD SUNPLL_SUNTR_PCHDL
xc1b Y YN net2 AVDD SUNPLL_SUNTR_PCHDL
xc2a net1 Y AVDD AVDD SUNPLL_SUNTR_PCHDL
xc2b YN Y net1 AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_ROSC <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_ROSC PWRUP_1V8 VDD_ROSC AVSS AVDD CK
xa3 N_2 N_1 CKUP CKDWN AVDD AVSS SUNPLL_SUN_PLL_LSCORE
xa40 CKUP CK AVDD AVSS SUNPLL_SUNTR_IVX1_CV
xa50 CKDWN NC1 AVDD AVSS SUNPLL_SUNTR_IVX1_CV
xa60 AVDD AVSS SUNPLL_SUNTR_TAPCELLB_CV
xb1 PWRUP_1V8 N_0 NI AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_NDX1_CV
xb2_0 NI N_7 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_1 N_7 N_6 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_2 N_6 N_5 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_3 N_5 N_4 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_4 N_4 N_3 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_5 N_3 N_2 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_6 N_2 N_1 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb2_7 N_1 N_0 AVDD AVSS VDD_ROSC AVSS SUNPLL_SUNTRB_IVX1_CV
xb3 AVDD AVSS SUNPLL_SUNTRB_TAPCELLBAVSS_CV
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_PFD <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_PFD CK_FB CK_REF CP_UP CP_DOWN AVDD AVSS
xa0 AVDD AVSS SUNPLL_SUNTR_TAPCELLB_CV
xa1 CFB CK_REF CP_UP_N AVDD AVSS SUNPLL_SUNTR_DFTSPCX1_CV
xa2 CP_UP_N CP_UP AVDD AVSS SUNPLL_SUNTR_IVX1_CV
xa3 CP_UP_N CP_DOWN_N CFB AVDD AVSS SUNPLL_SUNTR_NRX1_CV
xa5 CFB CK_FB CP_DOWN_N AVDD AVSS SUNPLL_SUNTR_DFTSPCX1_CV
xa6 CP_DOWN_N CP_DOWN AVDD AVSS SUNPLL_SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_DIVN <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_DIVN PWRUP_1V8 CK AVDD AVSS CK_FB
xa N0 D0 PWRUP_1V8 CK_FB N0 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
xb N1 D1 PWRUP_1V8 D0 N1 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
xc N2 D2 PWRUP_1V8 D1 N2 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
xd N3 D3 PWRUP_1V8 D2 N3 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
xe N4 D4 PWRUP_1V8 D3 N4 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
xf N5 D5 PWRUP_1V8 D4 N5 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
xg N6 CK PWRUP_1V8 D5 N6 AVDD AVSS SUNPLL_SUNTR_DFRNQNX1_CV
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_BUF <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_BUF AVDD VBN AVSS VI VO VFB
xa1 VS VBN AVSS AVSS SUNPLL_SUNTR_NCHDLCM
xa2 VDP VFB VS AVSS SUNPLL_SUNTR_NCHDLA
xa4 VGP VI VS AVSS SUNPLL_SUNTR_NCHDLA
xc1 VGP VDP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc2 VDP VDP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc3_0 VO VGP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc3_1 VO VGP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc3_2 VO VGP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc3_3 VO VGP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc3_4 VO VGP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xc3_5 VO VGP AVDD AVDD SUNPLL_SUNTR_PCHDLA
xd20 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd30 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd31 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd32 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd33 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd34 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd35 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd36 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd37 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xd38 VO AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_CP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_CP AVDD CP_UP_N CP_DOWN VBN AVSS LPF
xa10 VBP VBN AVSS AVSS SUNPLL_SUNTR_NCHDLCM
xa20 VNS VBN AVSS AVSS SUNPLL_SUNTR_NCHDLCM
xa30 LPF CP_DOWN VNS AVSS SUNPLL_SUNTR_NCHDL
xb10 VBP VBP AVDD AVDD SUNPLL_SUNTR_PCHDLCM
xb20 VPS VBP AVDD AVDD SUNPLL_SUNTR_PCHDLCM
xb30 LPF CP_UP_N VPS AVDD SUNPLL_SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_BIAS <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_BIAS IBPSR_1U AVDD PWRUP_1V8 AVSS
xa00 AVDD AVSS SUNPLL_SUNTR_TAPCELLB_CV
xa10 PWRUP_1V8 PWRUP_1V8_N AVDD AVSS SUNPLL_SUNTR_IVX1_CV
xa20 IBPSR_1U PWRUP_1V8_N AVSS AVSS SUNPLL_SUNTR_NCHDL
xa30 IBPSR_1U IBPSR_1U AVSS AVSS SUNPLL_SUNTR_NCHDLCM
.ENDS

*-------------------------------------------------------------
* SUNPLL_CAP_LPF <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_CAP_LPF A B
RR1 A NC0 sky130_fd_pr__res_generic_m1  l=0.4  w=0.4  
RR2 B NC1 sky130_fd_pr__res_generic_m1  l=0.4  w=0.4  
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL_LPF <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL_LPF VLPF AVSS
xa30 VN1 VLPF AVSS SUNPLL_SUNTR_RPPO_12k
xb10 VLPF AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb30 VLPF AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb31 VLPF AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb40 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb41 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb42 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb43 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb44 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb45 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb46 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb47 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb48 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
xb49 VN1 AVSS SUNPLL_SUNSAR_CAP_BSSW_CV
.ENDS

*-------------------------------------------------------------
* SUNPLL_SUN_PLL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNPLL_SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBSPR_1U
xb1 AVDD VDD_ROSC_N net2 VDD_ROSC_N IBSPR_1U AVSS SUNPLL_SUN_PLL_BUF
xb2 net2 AVSS SUNPLL_SUN_PLL_LPF
xh1 AVDD net1 CK PWRUP_1V8 AVSS SUNPLL_SUN_PLL_DIVN
xh2 AVDD CK VDD_ROSC_N PWRUP_1V8 AVSS SUNPLL_SUN_PLL_ROSC
xj1 AVDD CP_UP_N CK_REF CP_DOWN net1 AVSS SUNPLL_SUN_PLL_PFD
xk1 AVDD CP_UP_N net2 CP_DOWN IBSPR_1U AVSS SUNPLL_SUN_PLL_CP
xl2 IBSPR_1U AVDD PWRUP_1V8 AVSS SUNPLL_SUN_PLL_BIAS
.ENDS
