magic
tech sky130A
magscale 1 2
timestamp 1664582400
<< checkpaint >>
rect 0 0 5264 4236
<< locali >>
rect 16 16 5248 128
rect 16 16 5248 128
rect 16 16 128 4220
rect 16 4108 5248 4220
rect 5136 16 5248 4220
rect 16 16 5248 128
rect 4072 3438 4648 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 32 32 112 112
rect 112 32 192 112
rect 192 32 272 112
rect 272 32 352 112
rect 352 32 432 112
rect 432 32 512 112
rect 512 32 592 112
rect 592 32 672 112
rect 672 32 752 112
rect 752 32 832 112
rect 832 32 912 112
rect 912 32 992 112
rect 992 32 1072 112
rect 1072 32 1152 112
rect 1152 32 1232 112
rect 1232 32 1312 112
rect 1312 32 1392 112
rect 1392 32 1472 112
rect 1472 32 1552 112
rect 1552 32 1632 112
rect 1632 32 1712 112
rect 1712 32 1792 112
rect 1792 32 1872 112
rect 1872 32 1952 112
rect 1952 32 2032 112
rect 2032 32 2112 112
rect 2112 32 2192 112
rect 2192 32 2272 112
rect 2272 32 2352 112
rect 2352 32 2432 112
rect 2432 32 2512 112
rect 2512 32 2592 112
rect 2592 32 2672 112
rect 2672 32 2752 112
rect 2752 32 2832 112
rect 2832 32 2912 112
rect 2912 32 2992 112
rect 2992 32 3072 112
rect 3072 32 3152 112
rect 3152 32 3232 112
rect 3232 32 3312 112
rect 3312 32 3392 112
rect 3392 32 3472 112
rect 3472 32 3552 112
rect 3552 32 3632 112
rect 3632 32 3712 112
rect 3712 32 3792 112
rect 3792 32 3872 112
rect 3872 32 3952 112
rect 3952 32 4032 112
rect 4032 32 4112 112
rect 4112 32 4192 112
rect 4192 32 4272 112
rect 4272 32 4352 112
rect 4352 32 4432 112
rect 4432 32 4512 112
rect 4512 32 4592 112
rect 4592 32 4672 112
rect 4672 32 4752 112
rect 4752 32 4832 112
rect 4832 32 4912 112
rect 4912 32 4992 112
rect 4992 32 5072 112
rect 5072 32 5152 112
rect 5152 32 5232 112
rect 32 38 112 118
rect 32 118 112 198
rect 32 198 112 278
rect 32 278 112 358
rect 32 358 112 438
rect 32 438 112 518
rect 32 518 112 598
rect 32 598 112 678
rect 32 678 112 758
rect 32 758 112 838
rect 32 838 112 918
rect 32 918 112 998
rect 32 998 112 1078
rect 32 1078 112 1158
rect 32 1158 112 1238
rect 32 1238 112 1318
rect 32 1318 112 1398
rect 32 1398 112 1478
rect 32 1478 112 1558
rect 32 1558 112 1638
rect 32 1638 112 1718
rect 32 1718 112 1798
rect 32 1798 112 1878
rect 32 1878 112 1958
rect 32 1958 112 2038
rect 32 2038 112 2118
rect 32 2118 112 2198
rect 32 2198 112 2278
rect 32 2278 112 2358
rect 32 2358 112 2438
rect 32 2438 112 2518
rect 32 2518 112 2598
rect 32 2598 112 2678
rect 32 2678 112 2758
rect 32 2758 112 2838
rect 32 2838 112 2918
rect 32 2918 112 2998
rect 32 2998 112 3078
rect 32 3078 112 3158
rect 32 3158 112 3238
rect 32 3238 112 3318
rect 32 3318 112 3398
rect 32 3398 112 3478
rect 32 3478 112 3558
rect 32 3558 112 3638
rect 32 3638 112 3718
rect 32 3718 112 3798
rect 32 3798 112 3878
rect 32 3878 112 3958
rect 32 3958 112 4038
rect 32 4038 112 4118
rect 32 4118 112 4198
rect 32 4124 112 4204
rect 112 4124 192 4204
rect 192 4124 272 4204
rect 272 4124 352 4204
rect 352 4124 432 4204
rect 432 4124 512 4204
rect 512 4124 592 4204
rect 592 4124 672 4204
rect 672 4124 752 4204
rect 752 4124 832 4204
rect 832 4124 912 4204
rect 912 4124 992 4204
rect 992 4124 1072 4204
rect 1072 4124 1152 4204
rect 1152 4124 1232 4204
rect 1232 4124 1312 4204
rect 1312 4124 1392 4204
rect 1392 4124 1472 4204
rect 1472 4124 1552 4204
rect 1552 4124 1632 4204
rect 1632 4124 1712 4204
rect 1712 4124 1792 4204
rect 1792 4124 1872 4204
rect 1872 4124 1952 4204
rect 1952 4124 2032 4204
rect 2032 4124 2112 4204
rect 2112 4124 2192 4204
rect 2192 4124 2272 4204
rect 2272 4124 2352 4204
rect 2352 4124 2432 4204
rect 2432 4124 2512 4204
rect 2512 4124 2592 4204
rect 2592 4124 2672 4204
rect 2672 4124 2752 4204
rect 2752 4124 2832 4204
rect 2832 4124 2912 4204
rect 2912 4124 2992 4204
rect 2992 4124 3072 4204
rect 3072 4124 3152 4204
rect 3152 4124 3232 4204
rect 3232 4124 3312 4204
rect 3312 4124 3392 4204
rect 3392 4124 3472 4204
rect 3472 4124 3552 4204
rect 3552 4124 3632 4204
rect 3632 4124 3712 4204
rect 3712 4124 3792 4204
rect 3792 4124 3872 4204
rect 3872 4124 3952 4204
rect 3952 4124 4032 4204
rect 4032 4124 4112 4204
rect 4112 4124 4192 4204
rect 4192 4124 4272 4204
rect 4272 4124 4352 4204
rect 4352 4124 4432 4204
rect 4432 4124 4512 4204
rect 4512 4124 4592 4204
rect 4592 4124 4672 4204
rect 4672 4124 4752 4204
rect 4752 4124 4832 4204
rect 4832 4124 4912 4204
rect 4912 4124 4992 4204
rect 4992 4124 5072 4204
rect 5072 4124 5152 4204
rect 5152 4124 5232 4204
rect 5152 38 5232 118
rect 5152 118 5232 198
rect 5152 198 5232 278
rect 5152 278 5232 358
rect 5152 358 5232 438
rect 5152 438 5232 518
rect 5152 518 5232 598
rect 5152 598 5232 678
rect 5152 678 5232 758
rect 5152 758 5232 838
rect 5152 838 5232 918
rect 5152 918 5232 998
rect 5152 998 5232 1078
rect 5152 1078 5232 1158
rect 5152 1158 5232 1238
rect 5152 1238 5232 1318
rect 5152 1318 5232 1398
rect 5152 1398 5232 1478
rect 5152 1478 5232 1558
rect 5152 1558 5232 1638
rect 5152 1638 5232 1718
rect 5152 1718 5232 1798
rect 5152 1798 5232 1878
rect 5152 1878 5232 1958
rect 5152 1958 5232 2038
rect 5152 2038 5232 2118
rect 5152 2118 5232 2198
rect 5152 2198 5232 2278
rect 5152 2278 5232 2358
rect 5152 2358 5232 2438
rect 5152 2438 5232 2518
rect 5152 2518 5232 2598
rect 5152 2598 5232 2678
rect 5152 2678 5232 2758
rect 5152 2758 5232 2838
rect 5152 2838 5232 2918
rect 5152 2918 5232 2998
rect 5152 2998 5232 3078
rect 5152 3078 5232 3158
rect 5152 3158 5232 3238
rect 5152 3238 5232 3318
rect 5152 3318 5232 3398
rect 5152 3398 5232 3478
rect 5152 3478 5232 3558
rect 5152 3558 5232 3638
rect 5152 3638 5232 3718
rect 5152 3718 5232 3798
rect 5152 3798 5232 3878
rect 5152 3878 5232 3958
rect 5152 3958 5232 4038
rect 5152 4038 5232 4118
rect 5152 4118 5232 4198
<< ptap >>
rect 0 0 5264 144
rect 0 0 144 4236
rect 0 4092 5264 4236
rect 5120 0 5264 4236
use SUNTR_RES8 XA1
transform 1 0 688 0 1 688
box 688 688 4576 3548
<< labels >>
flabel locali s 16 16 5248 128 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 4072 3438 4648 3658 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
