magic
tech sky130A
magscale 1 2
timestamp 1660085871
<< checkpaint >>
rect -54 -592 11560 13728
<< m2 >>
rect 0 -592 11520 -288
rect 0 -592 11520 -288
rect 108 3190 334 3266
rect 334 836 1504 912
rect 334 1892 1504 1968
rect 334 2948 1504 3024
rect 334 836 410 3266
<< m3 >>
rect 6300 -592 6516 44
rect 6408 -44 11484 32
rect 6408 1012 11484 1088
rect 6408 2068 11484 2144
rect 6408 3124 11484 3200
rect 6408 4180 11484 4256
rect 6408 5236 11484 5312
rect 6408 6292 11484 6368
rect 6408 7348 11484 7424
rect 6408 8404 11484 8480
rect 6408 9460 11484 9536
rect 6408 10516 11484 10592
rect 6408 11572 11484 11648
rect 6408 12628 11484 12704
rect 11484 -44 11560 12704
<< locali >>
rect 216 -592 432 -88
rect -54 3190 270 3410
<< m1 >>
rect 540 3190 762 3250
rect 762 4004 1504 4064
rect 762 5060 1504 5120
rect 762 6116 1504 6176
rect 762 7172 1504 7232
rect 762 8228 1504 8288
rect 762 9284 1504 9344
rect 762 10340 1504 10400
rect 762 11396 1504 11456
rect 762 12452 1504 12512
rect 762 13508 1504 13568
rect 762 3190 822 13584
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_12k xa30
transform 1 0 0 0 1 440
box 0 440 648 3300
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb10
transform -1 0 11520 0 1 0
box 11520 0 21672 1056
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb30
transform -1 0 11520 0 1 1056
box 11520 1056 21672 2112
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb31
transform -1 0 11520 0 1 2112
box 11520 2112 21672 3168
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb40
transform -1 0 11520 0 1 3168
box 11520 3168 21672 4224
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb41
transform -1 0 11520 0 1 4224
box 11520 4224 21672 5280
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb42
transform -1 0 11520 0 1 5280
box 11520 5280 21672 6336
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb43
transform -1 0 11520 0 1 6336
box 11520 6336 21672 7392
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb44
transform -1 0 11520 0 1 7392
box 11520 7392 21672 8448
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb45
transform -1 0 11520 0 1 8448
box 11520 8448 21672 9504
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb46
transform -1 0 11520 0 1 9504
box 11520 9504 21672 10560
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb47
transform -1 0 11520 0 1 10560
box 11520 10560 21672 11616
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb48
transform -1 0 11520 0 1 11616
box 11520 11616 21672 12672
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xb49
transform -1 0 11520 0 1 12672
box 11520 12672 21672 13728
use cut_M3M4_2x1 
transform 1 0 6308 0 1 -592
box 6308 -592 6508 -516
use cut_M1M3_2x1 
transform 1 0 224 0 1 -592
box 224 -592 424 -516
use cut_M1M2_2x1 
transform 1 0 378 0 1 3190
box 378 3190 562 3258
use cut_M2M4_2x1 
transform 1 0 1404 0 1 4004
box 1404 4004 1604 4080
use cut_M2M4_2x1 
transform 1 0 1404 0 1 5060
box 1404 5060 1604 5136
use cut_M2M4_2x1 
transform 1 0 1404 0 1 6116
box 1404 6116 1604 6192
use cut_M2M4_2x1 
transform 1 0 1404 0 1 7172
box 1404 7172 1604 7248
use cut_M2M4_2x1 
transform 1 0 1404 0 1 8228
box 1404 8228 1604 8304
use cut_M2M4_2x1 
transform 1 0 1404 0 1 9284
box 1404 9284 1604 9360
use cut_M2M4_2x1 
transform 1 0 1404 0 1 10340
box 1404 10340 1604 10416
use cut_M2M4_2x1 
transform 1 0 1404 0 1 11396
box 1404 11396 1604 11472
use cut_M2M4_2x1 
transform 1 0 1404 0 1 12452
box 1404 12452 1604 12528
use cut_M2M4_2x1 
transform 1 0 1404 0 1 13508
box 1404 13508 1604 13584
use cut_M1M3_2x1 
transform 1 0 -54 0 1 3190
box -54 3190 146 3266
use cut_M3M4_2x1 
transform 1 0 1404 0 1 836
box 1404 836 1604 912
use cut_M3M4_2x1 
transform 1 0 1404 0 1 1892
box 1404 1892 1604 1968
use cut_M3M4_2x1 
transform 1 0 1404 0 1 2948
box 1404 2948 1604 3024
<< labels >>
flabel m2 s 0 -592 11520 -288 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s -54 3190 270 3410 0 FreeSans 400 0 0 0 VLPF
port 1 nsew
<< end >>
