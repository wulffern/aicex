magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 990 320
<< pdiff >>
rect 180 40 360 120
rect 180 120 360 200
rect 180 200 360 280
<< ntap >>
rect 900 -40 1080 40
rect 900 40 1080 120
rect 900 120 1080 200
rect 900 200 1080 280
rect 900 280 1080 360
<< poly >>
rect 120 -18 720 18
rect 120 142 720 178
rect 120 302 720 338
rect 540 120 720 200
<< pcontact >>
rect 560 140 600 160
rect 560 160 600 180
rect 600 140 660 160
rect 600 160 660 180
rect 660 140 700 160
rect 660 160 700 180
<< locali >>
rect 900 -40 1080 40
rect 180 50 360 110
rect 900 40 1080 120
rect 540 130 720 190
rect 900 120 1080 200
rect 180 210 360 270
rect 900 200 1080 280
rect 900 280 1080 360
<< ntapc >>
rect 960 40 1020 120
rect 960 120 1020 200
rect 960 200 1020 280
<< pdcontact >>
rect 200 60 240 80
rect 200 80 240 100
rect 240 60 300 80
rect 240 80 300 100
rect 300 60 340 80
rect 300 80 340 100
rect 200 220 240 240
rect 200 240 240 260
rect 240 220 300 240
rect 240 240 300 260
rect 300 220 340 240
rect 300 240 340 260
<< nwell >>
rect 0 -120 1140 440
<< labels >>
flabel locali s 540 130 720 190 0 FreeSans 400 0 0 0 G
port 1 nsew
flabel locali s 180 50 360 110 0 FreeSans 400 0 0 0 S
port 2 nsew
flabel locali s 900 120 1080 200 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 180 210 360 270 0 FreeSans 400 0 0 0 D
port 4 nsew
<< end >>
