magic
tech sky130A
magscale 1 2
timestamp 1658582973
<< checkpaint >>
rect -3928 -1848 28016 42182
<< m3 >>
rect 9100 18520 26178 18596
rect 9100 18908 26178 18984
rect 24104 19288 24180 26792
rect 24384 19288 24460 34536
rect 3944 19372 4020 30304
rect 4824 19566 4900 30304
rect 8984 19760 9060 30304
rect -216 19954 -140 30304
rect -216 19954 -140 30304
rect 13432 20148 13508 30330
rect 13432 20148 13508 30330
rect 18472 20342 18548 30330
rect 18472 20342 18548 30330
rect 10579 20536 10655 30330
rect 10579 20536 10655 30330
rect 15619 20730 15695 30330
rect 15619 20730 15695 30330
rect 499 20924 575 30330
rect 5539 21118 5615 30330
rect 5539 21118 5615 30330
rect 3352 21312 3428 30330
rect 3352 21312 3428 30330
rect 8392 21506 8468 30330
rect 8392 21506 8468 30330
rect 659 21700 735 31738
rect 8232 21894 8308 31738
rect 5699 22088 5775 31738
rect 3192 22282 3268 31738
rect 10914 22476 10990 33146
rect 13098 22670 13174 33146
rect 15954 22864 16030 33146
rect 8058 23058 8134 33146
rect 3018 23252 3094 33146
rect 834 23446 910 33146
rect 18138 23640 18214 33146
rect 5874 23834 5950 33146
rect 200 24534 400 40742
rect 3528 24534 3728 40742
rect 5240 24534 5440 40742
rect 8568 24534 8768 40742
rect 10280 24534 10480 40742
rect 13608 24534 13808 40742
rect 15320 24534 15520 40742
rect 18648 24534 18848 40742
rect 20360 24534 20560 40742
rect 23688 24534 23888 40742
rect 9648 -720 9848 5280
rect 14240 -720 14440 5280
rect 992 24534 1192 41462
rect 2736 24534 2936 41462
rect 6032 24534 6232 41462
rect 7776 24534 7976 41462
rect 11072 24534 11272 41462
rect 12816 24534 13016 41462
rect 16112 24534 16312 41462
rect 17856 24534 18056 41462
rect 21152 24534 21352 41462
rect 22896 24534 23096 41462
rect 8856 -1440 9056 5280
rect 15032 -1440 15232 5280
rect 1568 29344 1768 42182
rect 2160 29344 2360 42182
rect 6608 29344 6808 42182
rect 7200 29344 7400 42182
rect 11648 29344 11848 42182
rect 12240 29344 12440 42182
rect 16688 29344 16888 42182
rect 17280 29344 17480 42182
rect 21728 29344 21928 42182
rect 10294 -1848 10370 3470
rect 13718 -1848 13794 3470
rect 10924 1290 11180 1366
rect 9138 5474 10924 5550
rect 12908 1290 13088 1366
rect 13088 5474 14910 5550
rect 11180 1290 11360 1366
rect 11360 2698 12908 2774
rect 11360 1290 11436 2774
rect 11072 50 11272 126
rect 12816 50 13016 126
rect 20659 30330 20735 30530
<< m2 >>
rect 14872 18014 14948 18596
rect 9100 18014 9176 18984
rect 3944 19296 14020 19372
rect 4824 19490 13660 19566
rect 8984 19684 13300 19760
rect -216 19878 14380 19954
rect 11304 20072 13508 20148
rect 11664 20266 18548 20342
rect 10579 20460 11200 20536
rect 11484 20654 15695 20730
rect 499 20848 9760 20924
rect 5539 21042 10480 21118
rect 3352 21236 10120 21312
rect 8392 21430 10840 21506
rect 659 21624 9940 21700
rect 8232 21818 11020 21894
rect 5699 22012 10660 22088
rect 3192 22206 10300 22282
rect 10914 22400 12940 22476
rect 12684 22594 13174 22670
rect 12504 22788 16030 22864
rect 8058 22982 13120 23058
rect 3018 23176 13840 23252
rect 834 23370 14200 23446
rect 12324 23564 18214 23640
rect 5874 23758 13480 23834
rect 992 38526 1336 38602
rect 1336 37916 3944 37992
rect 3868 37916 3944 38116
rect 1336 37916 1412 38610
rect 6032 38526 6376 38602
rect 6376 37916 8984 37992
rect 8908 37916 8984 38116
rect 6376 37916 6452 38610
rect 11072 38526 11416 38602
rect 11416 37916 14024 37992
rect 13948 37916 14024 38116
rect 11416 37916 11492 38610
rect 16112 38526 16456 38602
rect 16456 37916 19064 37992
rect 18988 37916 19064 38116
rect 16456 37916 16532 38610
rect -232 34748 20144 34824
rect -308 34748 -232 34948
rect 3868 34748 3944 34948
rect 4732 34748 4808 34948
rect 8908 34748 8984 34948
rect 9772 34748 9848 34948
rect 13948 34748 14024 34948
rect 14812 34748 14888 34948
rect 18988 34748 19064 34948
rect 19852 34748 19928 34948
rect 1008 25288 1336 25364
rect 1336 24884 3944 24960
rect 3868 24884 3944 25100
rect 1336 24884 1412 25364
rect 6048 25288 6376 25364
rect 6376 24884 8984 24960
rect 8908 24884 8984 25100
rect 6376 24884 6452 25364
rect 11088 25288 11416 25364
rect 11416 24884 14024 24960
rect 13948 24884 14024 25100
rect 11416 24884 11492 25364
rect 16128 25288 16456 25364
rect 16456 24884 19064 24960
rect 18988 24884 19064 25100
rect 16456 24884 16532 25364
rect 21168 25288 21496 25364
rect 21496 25288 21572 25364
rect 2720 25288 3048 25364
rect 3048 25288 3124 25428
rect 3048 25428 4824 25504
rect 4748 25024 4824 25504
rect 7760 25288 8088 25364
rect 8088 25288 8164 25428
rect 8088 25428 9864 25504
rect 9788 25024 9864 25504
rect 12800 25288 13128 25364
rect 13128 25288 13204 25428
rect 13128 25428 14904 25504
rect 14828 25024 14904 25504
rect 17840 25288 18168 25364
rect 18168 25288 18244 25428
rect 18168 25428 19944 25504
rect 19868 25024 19944 25504
rect -216 27076 20144 27152
rect -292 26784 -216 27152
rect 3868 26784 3944 27152
rect 4748 26784 4824 27152
rect 8908 26784 8984 27152
rect 9788 26784 9864 27152
rect 13948 26784 14024 27152
rect 14828 26784 14904 27152
rect 18988 26784 19064 27152
rect 19868 26784 19944 27152
rect -232 27556 20144 27632
rect -308 27556 -232 27908
rect 3868 27556 3944 27908
rect 4732 27556 4808 27908
rect 8908 27556 8984 27908
rect 9772 27556 9848 27908
rect 13948 27556 14024 27908
rect 14812 27556 14888 27908
rect 18988 27556 19064 27908
rect 19852 27556 19928 27908
rect -16 28552 1424 28612
rect 1424 28552 1640 28612
rect 1424 28552 2504 28612
rect 1424 28552 6680 28612
rect 1424 28552 7544 28612
rect 1424 28552 11720 28612
rect 1424 28552 12584 28612
rect 1424 28552 16760 28612
rect 1424 28552 17624 28612
rect 1424 28552 21800 28612
rect 23396 30078 23780 30154
rect 20084 26860 23396 26936
rect 23396 26860 23472 30162
rect 20044 26784 20144 26860
rect 22740 31486 22988 31562
rect 20084 27924 22740 28000
rect 22740 27924 22816 31570
rect 20036 27848 20144 27924
rect 22556 38760 22728 38836
rect 20036 35592 22728 35668
rect 22728 35592 22804 38836
rect 22308 39464 22556 39540
rect 21260 38526 22308 38602
rect 22308 38526 22384 39540
rect 11180 2698 11352 2774
rect 11352 1290 12908 1366
rect 11352 1290 11428 2774
rect -232 28552 1640 28612
<< m4 >>
rect 24104 18908 24180 19288
rect 24384 18520 24460 19288
rect 10924 1290 11000 5550
rect 13088 1290 13164 5550
<< m1 >>
rect 13944 17954 14020 19296
rect 13584 17954 13660 19490
rect 13224 17954 13300 19684
rect 14304 17954 14380 19878
rect 11304 17954 11380 20072
rect 11664 17954 11740 20266
rect 11124 17954 11200 20460
rect 11484 17954 11560 20654
rect 9684 17954 9760 20848
rect 10404 17954 10480 21042
rect 10044 17954 10120 21236
rect 10764 17954 10840 21430
rect 9864 17954 9940 21624
rect 10944 17954 11020 21818
rect 10584 17954 10660 22012
rect 10224 17954 10300 22206
rect 12864 17954 12940 22400
rect 12684 17954 12760 22594
rect 12504 17954 12580 22788
rect 13044 17954 13120 22982
rect 13764 17954 13840 23176
rect 14124 17954 14200 23370
rect 12324 17954 12400 23564
rect 13404 17954 13480 23758
rect 10142 -1644 10202 558
rect 13886 -1644 13946 558
rect -3868 38056 -232 38116
rect 2720 38496 3056 38556
rect 3056 37936 4808 37996
rect 4748 37936 4808 38116
rect 3056 37936 3116 38564
rect 7760 38496 8096 38556
rect 8096 37936 9848 37996
rect 9788 37936 9848 38116
rect 8096 37936 8156 38564
rect 12800 38496 13136 38556
rect 13136 37936 14888 37996
rect 14828 37936 14888 38116
rect 13136 37936 13196 38564
rect 17840 38496 18176 38556
rect 18176 37936 19928 37996
rect 19868 37936 19928 38116
rect 18176 37936 18236 38564
rect 22328 39112 22556 39172
rect 20468 36384 22328 36444
rect 22328 36384 22388 39180
rect -3004 5474 76 5534
rect -3004 7034 76 7094
rect -3004 8594 76 8654
rect -3004 10154 76 10214
rect -3004 11714 76 11774
rect -3004 13274 76 13334
rect -3004 14834 76 14894
rect -3004 16394 76 16454
rect 23972 5474 27092 5534
rect 23972 7034 27092 7094
rect 23972 8594 27092 8654
rect 23972 10154 27092 10214
rect 23972 11714 27092 11774
rect 23972 13274 27092 13334
rect 23972 14834 27092 14894
rect 23972 16394 27092 16454
<< locali >>
rect 26892 -720 27092 40742
rect -3004 -720 27092 -520
rect -3004 40542 27092 40742
rect -3004 -720 -2804 40742
rect 26892 -720 27092 40742
rect 27612 -1440 27812 41462
rect -3724 -1440 27812 -1240
rect -3724 41262 27812 41462
rect -3724 -1440 -3524 41462
rect 27612 -1440 27812 41462
rect -3724 41982 27812 42182
rect -3724 41982 27812 42182
rect 27956 -1644 28016 42182
rect -3724 -1644 28016 -1584
rect 27956 -1644 28016 42182
rect -3928 -1848 28016 -1788
rect -3928 -1848 -3868 42182
rect 20360 36384 20576 36444
rect -232 34888 -16 34948
rect 1424 28552 1640 28612
rect 11072 2698 11288 2758
rect 11072 1290 11288 1350
use SARBSSW_CV XB1
transform -1 0 12044 0 1 0
box 12044 0 26372 5280
use SARBSSW_CV XB2
transform 1 0 12044 0 1 0
box 12044 0 26372 5280
use CDAC8_CV XDAC1
transform -1 0 11844 0 1 5474
box 11844 5474 23576 18014
use CDAC8_CV XDAC2
transform 1 0 12204 0 1 5474
box 12204 5474 23936 18014
use SARDIGEX4_CV XA0
transform 1 0 -556 0 1 24534
box -556 24534 1964 38966
use SARDIGEX4_CV XA1
transform -1 0 4484 0 1 24534
box 4484 24534 7004 38966
use SARDIGEX4_CV XA2
transform 1 0 4484 0 1 24534
box 4484 24534 7004 38966
use SARDIGEX4_CV XA3
transform -1 0 9524 0 1 24534
box 9524 24534 12044 38966
use SARDIGEX4_CV XA4
transform 1 0 9524 0 1 24534
box 9524 24534 12044 38966
use SARDIGEX4_CV XA5
transform -1 0 14564 0 1 24534
box 14564 24534 17084 38966
use SARDIGEX4_CV XA6
transform 1 0 14564 0 1 24534
box 14564 24534 17084 38966
use SARDIGEX4_CV XA7
transform -1 0 19604 0 1 24534
box 19604 24534 22124 38966
use SARDIGEX4_CV XA8
transform 1 0 19604 0 1 24534
box 19604 24534 22124 38966
use SARCMPX1_CV XA20
transform -1 0 24644 0 1 24534
box 24644 24534 27164 40022
use cut_M3M4_1x2 
transform 1 0 14872 0 1 18014
box 14872 18014 14948 18214
use cut_M3M4_2x1 
transform 1 0 14872 0 1 18520
box 14872 18520 15072 18596
use cut_M3M4_1x2 
transform 1 0 9100 0 1 18014
box 9100 18014 9176 18214
use cut_M3M4_2x1 
transform 1 0 9100 0 1 18908
box 9100 18908 9300 18984
use cut_M2M4_2x1 
transform 1 0 24104 0 1 26792
box 24104 26792 24304 26868
use cut_M4M5_2x1 
transform 1 0 24104 0 1 18908
box 24104 18908 24304 18984
use cut_M4M5_1x2 
transform 1 0 24104 0 1 19288
box 24104 19288 24180 19488
use cut_M3M4_2x1 
transform 1 0 24260 0 1 34536
box 24260 34536 24460 34612
use cut_M2M3_2x1 
transform 1 0 24104 0 1 34536
box 24104 34536 24304 34612
use cut_M4M5_2x1 
transform 1 0 24384 0 1 18520
box 24384 18520 24584 18596
use cut_M4M5_1x2 
transform 1 0 24384 0 1 19288
box 24384 19288 24460 19488
use cut_M3M4_1x2 
transform 1 0 3944 0 1 19234
box 3944 19234 4020 19434
use cut_M2M3_1x2 
transform 1 0 13936 0 1 19234
box 13936 19234 14012 19434
use cut_M3M4_1x2 
transform 1 0 4824 0 1 19428
box 4824 19428 4900 19628
use cut_M2M3_1x2 
transform 1 0 13576 0 1 19428
box 13576 19428 13652 19628
use cut_M3M4_1x2 
transform 1 0 8984 0 1 19622
box 8984 19622 9060 19822
use cut_M2M3_1x2 
transform 1 0 13216 0 1 19622
box 13216 19622 13292 19822
use cut_M3M4_1x2 
transform 1 0 -216 0 1 19816
box -216 19816 -140 20016
use cut_M2M3_1x2 
transform 1 0 14296 0 1 19816
box 14296 19816 14372 20016
use cut_M3M4_1x2 
transform 1 0 13432 0 1 20010
box 13432 20010 13508 20210
use cut_M2M3_1x2 
transform 1 0 11296 0 1 20010
box 11296 20010 11372 20210
use cut_M3M4_1x2 
transform 1 0 18472 0 1 20204
box 18472 20204 18548 20404
use cut_M2M3_1x2 
transform 1 0 11656 0 1 20204
box 11656 20204 11732 20404
use cut_M3M4_1x2 
transform 1 0 10579 0 1 20398
box 10579 20398 10655 20598
use cut_M2M3_1x2 
transform 1 0 11116 0 1 20398
box 11116 20398 11192 20598
use cut_M3M4_1x2 
transform 1 0 15619 0 1 20592
box 15619 20592 15695 20792
use cut_M2M3_1x2 
transform 1 0 11476 0 1 20592
box 11476 20592 11552 20792
use cut_M3M4_1x2 
transform 1 0 499 0 1 20786
box 499 20786 575 20986
use cut_M2M3_1x2 
transform 1 0 9676 0 1 20786
box 9676 20786 9752 20986
use cut_M3M4_1x2 
transform 1 0 5539 0 1 20980
box 5539 20980 5615 21180
use cut_M2M3_1x2 
transform 1 0 10396 0 1 20980
box 10396 20980 10472 21180
use cut_M3M4_1x2 
transform 1 0 3352 0 1 21174
box 3352 21174 3428 21374
use cut_M2M3_1x2 
transform 1 0 10036 0 1 21174
box 10036 21174 10112 21374
use cut_M3M4_1x2 
transform 1 0 8392 0 1 21368
box 8392 21368 8468 21568
use cut_M2M3_1x2 
transform 1 0 10756 0 1 21368
box 10756 21368 10832 21568
use cut_M3M4_1x2 
transform 1 0 659 0 1 21562
box 659 21562 735 21762
use cut_M2M3_1x2 
transform 1 0 9856 0 1 21562
box 9856 21562 9932 21762
use cut_M3M4_1x2 
transform 1 0 8232 0 1 21756
box 8232 21756 8308 21956
use cut_M2M3_1x2 
transform 1 0 10936 0 1 21756
box 10936 21756 11012 21956
use cut_M3M4_1x2 
transform 1 0 5699 0 1 21950
box 5699 21950 5775 22150
use cut_M2M3_1x2 
transform 1 0 10576 0 1 21950
box 10576 21950 10652 22150
use cut_M3M4_1x2 
transform 1 0 3192 0 1 22144
box 3192 22144 3268 22344
use cut_M2M3_1x2 
transform 1 0 10216 0 1 22144
box 10216 22144 10292 22344
use cut_M3M4_1x2 
transform 1 0 10914 0 1 22338
box 10914 22338 10990 22538
use cut_M2M3_1x2 
transform 1 0 12856 0 1 22338
box 12856 22338 12932 22538
use cut_M3M4_1x2 
transform 1 0 13098 0 1 22532
box 13098 22532 13174 22732
use cut_M2M3_1x2 
transform 1 0 12676 0 1 22532
box 12676 22532 12752 22732
use cut_M3M4_1x2 
transform 1 0 15954 0 1 22726
box 15954 22726 16030 22926
use cut_M2M3_1x2 
transform 1 0 12496 0 1 22726
box 12496 22726 12572 22926
use cut_M3M4_1x2 
transform 1 0 8058 0 1 22920
box 8058 22920 8134 23120
use cut_M2M3_1x2 
transform 1 0 13036 0 1 22920
box 13036 22920 13112 23120
use cut_M3M4_1x2 
transform 1 0 3018 0 1 23114
box 3018 23114 3094 23314
use cut_M2M3_1x2 
transform 1 0 13756 0 1 23114
box 13756 23114 13832 23314
use cut_M3M4_1x2 
transform 1 0 834 0 1 23308
box 834 23308 910 23508
use cut_M2M3_1x2 
transform 1 0 14116 0 1 23308
box 14116 23308 14192 23508
use cut_M3M4_1x2 
transform 1 0 18138 0 1 23502
box 18138 23502 18214 23702
use cut_M2M3_1x2 
transform 1 0 12316 0 1 23502
box 12316 23502 12392 23702
use cut_M3M4_1x2 
transform 1 0 5874 0 1 23696
box 5874 23696 5950 23896
use cut_M2M3_1x2 
transform 1 0 13396 0 1 23696
box 13396 23696 13472 23896
use cut_M1M4_2x2 
transform 1 0 200 0 1 40542
box 200 40542 400 40742
use cut_M1M4_2x2 
transform 1 0 3528 0 1 40542
box 3528 40542 3728 40742
use cut_M1M4_2x2 
transform 1 0 5240 0 1 40542
box 5240 40542 5440 40742
use cut_M1M4_2x2 
transform 1 0 8568 0 1 40542
box 8568 40542 8768 40742
use cut_M1M4_2x2 
transform 1 0 10280 0 1 40542
box 10280 40542 10480 40742
use cut_M1M4_2x2 
transform 1 0 13608 0 1 40542
box 13608 40542 13808 40742
use cut_M1M4_2x2 
transform 1 0 15320 0 1 40542
box 15320 40542 15520 40742
use cut_M1M4_2x2 
transform 1 0 18648 0 1 40542
box 18648 40542 18848 40742
use cut_M1M4_2x2 
transform 1 0 20360 0 1 40542
box 20360 40542 20560 40742
use cut_M1M4_2x2 
transform 1 0 23688 0 1 40542
box 23688 40542 23888 40742
use cut_M1M4_2x2 
transform 1 0 9648 0 1 -720
box 9648 -720 9848 -520
use cut_M1M4_2x2 
transform 1 0 14240 0 1 -720
box 14240 -720 14440 -520
use cut_M1M4_2x2 
transform 1 0 992 0 1 41262
box 992 41262 1192 41462
use cut_M1M4_2x2 
transform 1 0 2736 0 1 41262
box 2736 41262 2936 41462
use cut_M1M4_2x2 
transform 1 0 6032 0 1 41262
box 6032 41262 6232 41462
use cut_M1M4_2x2 
transform 1 0 7776 0 1 41262
box 7776 41262 7976 41462
use cut_M1M4_2x2 
transform 1 0 11072 0 1 41262
box 11072 41262 11272 41462
use cut_M1M4_2x2 
transform 1 0 12816 0 1 41262
box 12816 41262 13016 41462
use cut_M1M4_2x2 
transform 1 0 16112 0 1 41262
box 16112 41262 16312 41462
use cut_M1M4_2x2 
transform 1 0 17856 0 1 41262
box 17856 41262 18056 41462
use cut_M1M4_2x2 
transform 1 0 21152 0 1 41262
box 21152 41262 21352 41462
use cut_M1M4_2x2 
transform 1 0 22896 0 1 41262
box 22896 41262 23096 41462
use cut_M1M4_2x2 
transform 1 0 8856 0 1 -1440
box 8856 -1440 9056 -1240
use cut_M1M4_2x2 
transform 1 0 15032 0 1 -1440
box 15032 -1440 15232 -1240
use cut_M1M4_2x2 
transform 1 0 1568 0 1 41982
box 1568 41982 1768 42182
use cut_M1M4_2x2 
transform 1 0 2160 0 1 41982
box 2160 41982 2360 42182
use cut_M1M4_2x2 
transform 1 0 6608 0 1 41982
box 6608 41982 6808 42182
use cut_M1M4_2x2 
transform 1 0 7200 0 1 41982
box 7200 41982 7400 42182
use cut_M1M4_2x2 
transform 1 0 11648 0 1 41982
box 11648 41982 11848 42182
use cut_M1M4_2x2 
transform 1 0 12240 0 1 41982
box 12240 41982 12440 42182
use cut_M1M4_2x2 
transform 1 0 16688 0 1 41982
box 16688 41982 16888 42182
use cut_M1M4_2x2 
transform 1 0 17280 0 1 41982
box 17280 41982 17480 42182
use cut_M1M4_2x2 
transform 1 0 21728 0 1 41982
box 21728 41982 21928 42182
use cut_M1M2_2x1 
transform 1 0 10080 0 1 498
box 10080 498 10264 566
use cut_M1M2_2x1 
transform 1 0 10080 0 1 -1644
box 10080 -1644 10264 -1576
use cut_M1M2_2x1 
transform 1 0 13824 0 1 498
box 13824 498 14008 566
use cut_M1M2_2x1 
transform 1 0 13824 0 1 -1644
box 13824 -1644 14008 -1576
use cut_M1M2_2x1 
transform 1 0 -232 0 1 38056
box -232 38056 -48 38124
use cut_M1M2_1x2 
transform 1 0 -3932 0 1 37994
box -3932 37994 -3864 38178
use cut_M1M4_2x1 
transform 1 0 10232 0 1 -1848
box 10232 -1848 10432 -1772
use cut_M1M4_2x1 
transform 1 0 13656 0 1 -1848
box 13656 -1848 13856 -1772
use cut_M1M3_2x1 
transform 1 0 992 0 1 38534
box 992 38534 1192 38610
use cut_M1M3_2x1 
transform 1 0 3944 0 1 38056
box 3944 38056 4144 38132
use cut_M1M3_2x1 
transform 1 0 6032 0 1 38534
box 6032 38534 6232 38610
use cut_M1M3_2x1 
transform 1 0 8984 0 1 38056
box 8984 38056 9184 38132
use cut_M1M3_2x1 
transform 1 0 11072 0 1 38534
box 11072 38534 11272 38610
use cut_M1M3_2x1 
transform 1 0 14024 0 1 38056
box 14024 38056 14224 38132
use cut_M1M3_2x1 
transform 1 0 16112 0 1 38534
box 16112 38534 16312 38610
use cut_M1M3_2x1 
transform 1 0 19064 0 1 38056
box 19064 38056 19264 38132
use cut_M1M3_2x1 
transform 1 0 -232 0 1 34888
box -232 34888 -32 34964
use cut_M1M3_2x1 
transform 1 0 3944 0 1 34888
box 3944 34888 4144 34964
use cut_M1M3_2x1 
transform 1 0 4808 0 1 34888
box 4808 34888 5008 34964
use cut_M1M3_2x1 
transform 1 0 8984 0 1 34888
box 8984 34888 9184 34964
use cut_M1M3_2x1 
transform 1 0 9848 0 1 34888
box 9848 34888 10048 34964
use cut_M1M3_2x1 
transform 1 0 14024 0 1 34888
box 14024 34888 14224 34964
use cut_M1M3_2x1 
transform 1 0 14888 0 1 34888
box 14888 34888 15088 34964
use cut_M1M3_2x1 
transform 1 0 19064 0 1 34888
box 19064 34888 19264 34964
use cut_M1M3_2x1 
transform 1 0 19928 0 1 34888
box 19928 34888 20128 34964
use cut_M1M2_2x1 
transform 1 0 2720 0 1 38496
box 2720 38496 2904 38564
use cut_M1M2_2x1 
transform 1 0 4808 0 1 38056
box 4808 38056 4992 38124
use cut_M1M2_2x1 
transform 1 0 7760 0 1 38496
box 7760 38496 7944 38564
use cut_M1M2_2x1 
transform 1 0 9848 0 1 38056
box 9848 38056 10032 38124
use cut_M1M2_2x1 
transform 1 0 12800 0 1 38496
box 12800 38496 12984 38564
use cut_M1M2_2x1 
transform 1 0 14888 0 1 38056
box 14888 38056 15072 38124
use cut_M1M2_2x1 
transform 1 0 17840 0 1 38496
box 17840 38496 18024 38564
use cut_M1M2_2x1 
transform 1 0 19928 0 1 38056
box 19928 38056 20112 38124
use cut_M1M3_2x1 
transform 1 0 -232 0 1 27848
box -232 27848 -32 27924
use cut_M1M3_2x1 
transform 1 0 3944 0 1 27848
box 3944 27848 4144 27924
use cut_M1M3_2x1 
transform 1 0 4808 0 1 27848
box 4808 27848 5008 27924
use cut_M1M3_2x1 
transform 1 0 8984 0 1 27848
box 8984 27848 9184 27924
use cut_M1M3_2x1 
transform 1 0 9848 0 1 27848
box 9848 27848 10048 27924
use cut_M1M3_2x1 
transform 1 0 14024 0 1 27848
box 14024 27848 14224 27924
use cut_M1M3_2x1 
transform 1 0 14888 0 1 27848
box 14888 27848 15088 27924
use cut_M1M3_2x1 
transform 1 0 19064 0 1 27848
box 19064 27848 19264 27924
use cut_M1M3_2x1 
transform 1 0 19928 0 1 27848
box 19928 27848 20128 27924
use cut_M1M3_2x1 
transform 1 0 1424 0 1 28552
box 1424 28552 1624 28628
use cut_M1M3_2x1 
transform 1 0 1424 0 1 28552
box 1424 28552 1624 28628
use cut_M1M3_2x1 
transform 1 0 2288 0 1 28552
box 2288 28552 2488 28628
use cut_M1M3_2x1 
transform 1 0 6464 0 1 28552
box 6464 28552 6664 28628
use cut_M1M3_2x1 
transform 1 0 7328 0 1 28552
box 7328 28552 7528 28628
use cut_M1M3_2x1 
transform 1 0 11504 0 1 28552
box 11504 28552 11704 28628
use cut_M1M3_2x1 
transform 1 0 12368 0 1 28552
box 12368 28552 12568 28628
use cut_M1M3_2x1 
transform 1 0 16544 0 1 28552
box 16544 28552 16744 28628
use cut_M1M3_2x1 
transform 1 0 17408 0 1 28552
box 17408 28552 17608 28628
use cut_M1M3_2x1 
transform 1 0 21584 0 1 28552
box 21584 28552 21784 28628
use cut_M1M3_2x1 
transform 1 0 23688 0 1 30086
box 23688 30086 23888 30162
use cut_M1M3_2x1 
transform 1 0 22896 0 1 31494
box 22896 31494 23096 31570
use cut_M1M3_2x1 
transform 1 0 22448 0 1 38760
box 22448 38760 22648 38836
use cut_M1M3_2x1 
transform 1 0 19928 0 1 35592
box 19928 35592 20128 35668
use cut_M1M3_2x1 
transform 1 0 22464 0 1 39464
box 22464 39464 22664 39540
use cut_M1M3_2x1 
transform 1 0 21168 0 1 38534
box 21168 38534 21368 38610
use cut_M1M2_2x1 
transform 1 0 22480 0 1 39112
box 22480 39112 22664 39180
use cut_M1M2_2x1 
transform 1 0 20392 0 1 36384
box 20392 36384 20576 36452
use cut_M4M5_1x2 
transform 1 0 10924 0 1 1290
box 10924 1290 11000 1490
use cut_M4M5_1x2 
transform 1 0 10924 0 1 5350
box 10924 5350 11000 5550
use cut_M1M4_2x1 
transform 1 0 12800 0 1 1290
box 12800 1290 13000 1366
use cut_M4M5_1x2 
transform 1 0 13088 0 1 1290
box 13088 1290 13164 1490
use cut_M4M5_1x2 
transform 1 0 13088 0 1 5350
box 13088 5350 13164 5550
use cut_M1M3_2x1 
transform 1 0 11072 0 1 2698
box 11072 2698 11272 2774
use cut_M1M3_2x1 
transform 1 0 12800 0 1 1290
box 12800 1290 13000 1366
use cut_M1M4_2x1 
transform 1 0 11072 0 1 1290
box 11072 1290 11272 1366
use cut_M1M4_2x1 
transform 1 0 12800 0 1 2698
box 12800 2698 13000 2774
use cut_M1M3_2x1 
transform 1 0 -232 0 1 28552
box -232 28552 -32 28628
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 5534
box -3004 5534 -2820 5718
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 7094
box -3004 7094 -2820 7278
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 8654
box -3004 8654 -2820 8838
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 10214
box -3004 10214 -2820 10398
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 11774
box -3004 11774 -2820 11958
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 13334
box -3004 13334 -2820 13518
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 14894
box -3004 14894 -2820 15078
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 16454
box -3004 16454 -2820 16638
use cut_M1M2_2x2 
transform 1 0 26908 0 1 5474
box 26908 5474 27092 5658
use cut_M1M2_2x2 
transform 1 0 26908 0 1 7034
box 26908 7034 27092 7218
use cut_M1M2_2x2 
transform 1 0 26908 0 1 8594
box 26908 8594 27092 8778
use cut_M1M2_2x2 
transform 1 0 26908 0 1 10154
box 26908 10154 27092 10338
use cut_M1M2_2x2 
transform 1 0 26908 0 1 11714
box 26908 11714 27092 11898
use cut_M1M2_2x2 
transform 1 0 26908 0 1 13274
box 26908 13274 27092 13458
use cut_M1M2_2x2 
transform 1 0 26908 0 1 14834
box 26908 14834 27092 15018
use cut_M1M2_2x2 
transform 1 0 26908 0 1 16394
box 26908 16394 27092 16578
<< labels >>
flabel m3 s -216 19954 -140 30304 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 13432 20148 13508 30330 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 18472 20342 18548 30330 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 10579 20536 10655 30330 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 15619 20730 15695 30330 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 5539 21118 5615 30330 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 3352 21312 3428 30330 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8392 21506 8468 30330 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel locali s 26892 -720 27092 40742 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
flabel locali s 27612 -1440 27812 41462 0 FreeSans 400 0 0 0 AVDD
port 10 nsew
flabel locali s -3724 41982 27812 42182 0 FreeSans 400 0 0 0 VREF
port 11 nsew
flabel locali s 27956 -1644 28016 42182 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 12 nsew
flabel locali s 20360 36384 20576 36444 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 11072 50 11272 126 0 FreeSans 400 0 0 0 SAR_IP
port 14 nsew
flabel m3 s 12816 50 13016 126 0 FreeSans 400 0 0 0 SAR_IN
port 15 nsew
flabel locali s -232 34888 -16 34948 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 1424 28552 1640 28612 0 FreeSans 400 0 0 0 EN
port 17 nsew
flabel locali s 11072 2698 11288 2758 0 FreeSans 400 0 0 0 SARN
port 18 nsew
flabel locali s 11072 1290 11288 1350 0 FreeSans 400 0 0 0 SARP
port 19 nsew
flabel m3 s 20659 30330 20735 30530 0 FreeSans 400 0 0 0 D<0>
port 20 nsew
<< end >>
