magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 30 8960 1518
<< m3 >>
rect 312 0 380 1548
rect 312 0 380 1548
rect 444 132 512 1416
rect 576 0 644 1548
rect 708 132 776 1416
rect 840 0 908 1548
rect 972 132 1040 1416
rect 1104 0 1172 1548
rect 1236 132 1304 1416
rect 1368 0 1436 1548
rect 1500 132 1568 1416
rect 1632 0 1700 1548
rect 1764 132 1832 1416
rect 1896 0 1964 1548
rect 2028 132 2096 1416
rect 2160 0 2228 1548
rect 2292 132 2360 1416
rect 2424 0 2492 1548
rect 2556 132 2624 1416
rect 2688 0 2756 1548
rect 2820 132 2888 1416
rect 2952 0 3020 1548
rect 3084 132 3152 1416
rect 3216 0 3284 1548
rect 3348 132 3416 1416
rect 3480 0 3548 1548
rect 3612 132 3680 1416
rect 3744 0 3812 1548
rect 3876 132 3944 1416
rect 4008 0 4076 1548
rect 4140 132 4208 1416
rect 4272 0 4340 1548
rect 4404 132 4472 1416
rect 4536 0 4604 1548
rect 4668 132 4736 1416
rect 4800 0 4868 1548
rect 4932 132 5000 1416
rect 5064 0 5132 1548
rect 5196 132 5264 1416
rect 5328 0 5396 1548
rect 5460 132 5528 1416
rect 5592 0 5660 1548
rect 5724 132 5792 1416
rect 5856 0 5924 1548
rect 5988 132 6056 1416
rect 6120 0 6188 1548
rect 6252 132 6320 1416
rect 6384 0 6452 1548
rect 6516 132 6584 1416
rect 6648 0 6716 1548
rect 6780 132 6848 1416
rect 6912 0 6980 1548
rect 7044 132 7112 1416
rect 7176 0 7244 1548
rect 7308 132 7376 1416
rect 7440 0 7508 1548
rect 7572 132 7640 1416
rect 7704 0 7772 1548
rect 7836 132 7904 1416
rect 7968 0 8036 1548
rect 8100 132 8168 1416
rect 8232 0 8300 1548
rect 8364 132 8432 1416
rect 8496 0 8564 1548
rect 8628 132 8696 1416
rect 8892 0 8960 1548
rect 8760 0 8828 1548
rect 312 0 8760 68
rect 312 1480 8760 1548
<< m1 >>
rect 312 0 8892 68
rect 2292 380 2360 1548
rect 6780 0 6848 1168
rect 2556 0 2624 508
rect 2556 820 2624 1548
rect 6516 0 6584 508
rect 6516 820 6584 1548
rect 2028 0 2096 948
rect 2028 1260 2096 1548
rect 2820 0 2888 948
rect 2820 1260 2888 1548
rect 6252 0 6320 948
rect 6252 1260 6320 1548
rect 7044 0 7112 948
rect 7044 1260 7112 1548
rect 1500 0 1568 728
rect 1500 1040 1568 1548
rect 1764 0 1832 728
rect 1764 1040 1832 1548
rect 3084 0 3152 728
rect 3084 1040 3152 1548
rect 3348 0 3416 728
rect 3348 1040 3416 1548
rect 5724 0 5792 728
rect 5724 1040 5792 1548
rect 5988 0 6056 728
rect 5988 1040 6056 1548
rect 7308 0 7376 728
rect 7308 1040 7376 1548
rect 7572 0 7640 728
rect 7572 1040 7640 1548
rect 444 0 512 288
rect 444 600 512 1548
rect 708 0 776 288
rect 708 600 776 1548
rect 972 0 1040 288
rect 972 600 1040 1548
rect 1236 0 1304 288
rect 1236 600 1304 1548
rect 3612 0 3680 288
rect 3612 600 3680 1548
rect 3876 0 3944 288
rect 3876 600 3944 1548
rect 4140 0 4208 288
rect 4140 600 4208 1548
rect 4404 0 4472 288
rect 4404 600 4472 1548
rect 4668 0 4736 288
rect 4668 600 4736 1548
rect 4932 0 5000 288
rect 4932 600 5000 1548
rect 5196 0 5264 288
rect 5196 600 5264 1548
rect 5460 0 5528 288
rect 5460 600 5528 1548
rect 7836 0 7904 288
rect 7836 600 7904 1548
rect 8100 0 8168 288
rect 8100 600 8168 1548
rect 8364 0 8432 288
rect 8364 600 8432 1548
rect 8628 0 8696 288
rect 8628 600 8696 1548
rect 312 0 380 1480
rect 576 0 644 1480
rect 840 0 908 1480
rect 1104 0 1172 1480
rect 1368 0 1436 1480
rect 1632 0 1700 1480
rect 1896 0 1964 1480
rect 2160 0 2228 1480
rect 2424 0 2492 1480
rect 2688 0 2756 1480
rect 2952 0 3020 1480
rect 3216 0 3284 1480
rect 3480 0 3548 1480
rect 3744 0 3812 1480
rect 4008 0 4076 1480
rect 4272 0 4340 1480
rect 4536 0 4604 1480
rect 4800 0 4868 1480
rect 5064 0 5132 1480
rect 5328 0 5396 1480
rect 5592 0 5660 1480
rect 5856 0 5924 1480
rect 6120 0 6188 1480
rect 6384 0 6452 1480
rect 6648 0 6716 1480
rect 6912 0 6980 1480
rect 7176 0 7244 1480
rect 7440 0 7508 1480
rect 7704 0 7772 1480
rect 7968 0 8036 1480
rect 8232 0 8300 1480
rect 8496 0 8564 1480
rect 8892 0 8960 1548
rect 8760 0 8828 1548
rect 312 0 8892 68
rect 312 1480 8892 1548
<< locali >>
rect 0 190 184 258
rect 0 1290 184 1358
rect 0 630 184 698
rect 0 1070 184 1138
rect 0 850 184 918
rect 0 410 184 478
rect 0 410 8760 478
rect 0 190 8760 258
rect 0 1290 8760 1358
rect 0 630 8760 698
rect 0 1070 8760 1138
rect 0 850 8760 918
<< m4 >>
rect 180 0 248 1548
rect 444 0 512 1548
rect 708 0 776 1548
rect 972 0 1040 1548
rect 1236 0 1304 1548
rect 1500 0 1568 1548
rect 1764 0 1832 1548
rect 2028 0 2096 1548
rect 2292 0 2360 1548
rect 2556 0 2624 1548
rect 2820 0 2888 1548
rect 3084 0 3152 1548
rect 3348 0 3416 1548
rect 3612 0 3680 1548
rect 3876 0 3944 1548
rect 4140 0 4208 1548
rect 4404 0 4472 1548
rect 4668 0 4736 1548
rect 4932 0 5000 1548
rect 5196 0 5264 1548
rect 5460 0 5528 1548
rect 5724 0 5792 1548
rect 5988 0 6056 1548
rect 6252 0 6320 1548
rect 6516 0 6584 1548
rect 6780 0 6848 1548
rect 7044 0 7112 1548
rect 7308 0 7376 1548
rect 7572 0 7640 1548
rect 7836 0 7904 1548
rect 8100 0 8168 1548
rect 8364 0 8432 1548
rect 8628 0 8696 1548
rect 8892 0 8960 1548
rect 180 0 8892 68
rect 180 1480 8892 1548
<< m2 >>
rect 444 132 512 1416
rect 708 132 776 1416
rect 972 132 1040 1416
rect 1236 132 1304 1416
rect 1500 132 1568 1416
rect 1764 132 1832 1416
rect 2028 132 2096 1416
rect 2292 132 2360 1416
rect 2556 132 2624 1416
rect 2820 132 2888 1416
rect 3084 132 3152 1416
rect 3348 132 3416 1416
rect 3612 132 3680 1416
rect 3876 132 3944 1416
rect 4140 132 4208 1416
rect 4404 132 4472 1416
rect 4668 132 4736 1416
rect 4932 132 5000 1416
rect 5196 132 5264 1416
rect 5460 132 5528 1416
rect 5724 132 5792 1416
rect 5988 132 6056 1416
rect 6252 132 6320 1416
rect 6516 132 6584 1416
rect 6780 132 6848 1416
rect 7044 132 7112 1416
rect 7308 132 7376 1416
rect 7572 132 7640 1416
rect 7836 132 7904 1416
rect 8100 132 8168 1416
rect 8364 132 8432 1416
rect 8628 132 8696 1416
rect 8892 0 8960 1548
use RM1 XRES1A
transform 1 0 184 0 1 190
box 184 190 304 190
use RM1 XRES1B
transform 1 0 184 0 1 1290
box 184 1290 304 1290
use RM1 XRES2
transform 1 0 184 0 1 630
box 184 630 304 630
use RM1 XRES4
transform 1 0 184 0 1 1070
box 184 1070 304 1070
use RM1 XRES8
transform 1 0 184 0 1 850
box 184 850 304 850
use RM1 XRES16
transform 1 0 184 0 1 410
box 184 410 304 410
use cut_M2M5_1x2 
transform 1 0 8892 0 1 590
box 8892 590 8960 774
use cut_M1M4_1x2 
transform 1 0 2292 0 1 132
box 2292 132 2360 316
use cut_M1M4_1x2 
transform 1 0 6780 0 1 1232
box 6780 1232 6848 1416
use cut_M1M4_1x2 
transform 1 0 2556 0 1 572
box 2556 572 2624 756
use cut_M1M4_1x2 
transform 1 0 6516 0 1 572
box 6516 572 6584 756
use cut_M1M4_1x2 
transform 1 0 2028 0 1 1012
box 2028 1012 2096 1196
use cut_M1M4_1x2 
transform 1 0 2820 0 1 1012
box 2820 1012 2888 1196
use cut_M1M4_1x2 
transform 1 0 6252 0 1 1012
box 6252 1012 6320 1196
use cut_M1M4_1x2 
transform 1 0 7044 0 1 1012
box 7044 1012 7112 1196
use cut_M1M4_1x2 
transform 1 0 1500 0 1 792
box 1500 792 1568 976
use cut_M1M4_1x2 
transform 1 0 1764 0 1 792
box 1764 792 1832 976
use cut_M1M4_1x2 
transform 1 0 3084 0 1 792
box 3084 792 3152 976
use cut_M1M4_1x2 
transform 1 0 3348 0 1 792
box 3348 792 3416 976
use cut_M1M4_1x2 
transform 1 0 5724 0 1 792
box 5724 792 5792 976
use cut_M1M4_1x2 
transform 1 0 5988 0 1 792
box 5988 792 6056 976
use cut_M1M4_1x2 
transform 1 0 7308 0 1 792
box 7308 792 7376 976
use cut_M1M4_1x2 
transform 1 0 7572 0 1 792
box 7572 792 7640 976
use cut_M1M4_1x2 
transform 1 0 444 0 1 352
box 444 352 512 536
use cut_M1M4_1x2 
transform 1 0 708 0 1 352
box 708 352 776 536
use cut_M1M4_1x2 
transform 1 0 972 0 1 352
box 972 352 1040 536
use cut_M1M4_1x2 
transform 1 0 1236 0 1 352
box 1236 352 1304 536
use cut_M1M4_1x2 
transform 1 0 3612 0 1 352
box 3612 352 3680 536
use cut_M1M4_1x2 
transform 1 0 3876 0 1 352
box 3876 352 3944 536
use cut_M1M4_1x2 
transform 1 0 4140 0 1 352
box 4140 352 4208 536
use cut_M1M4_1x2 
transform 1 0 4404 0 1 352
box 4404 352 4472 536
use cut_M1M4_1x2 
transform 1 0 4668 0 1 352
box 4668 352 4736 536
use cut_M1M4_1x2 
transform 1 0 4932 0 1 352
box 4932 352 5000 536
use cut_M1M4_1x2 
transform 1 0 5196 0 1 352
box 5196 352 5264 536
use cut_M1M4_1x2 
transform 1 0 5460 0 1 352
box 5460 352 5528 536
use cut_M1M4_1x2 
transform 1 0 7836 0 1 352
box 7836 352 7904 536
use cut_M1M4_1x2 
transform 1 0 8100 0 1 352
box 8100 352 8168 536
use cut_M1M4_1x2 
transform 1 0 8364 0 1 352
box 8364 352 8432 536
use cut_M1M4_1x2 
transform 1 0 8628 0 1 352
box 8628 352 8696 536
<< labels >>
flabel m3 s 312 0 380 1548 0 FreeSans 400 0 0 0 CTOP
port 1 nsew
flabel m1 s 312 0 8892 68 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 0 190 184 258 0 FreeSans 400 0 0 0 C1A
port 3 nsew
flabel locali s 0 1290 184 1358 0 FreeSans 400 0 0 0 C1B
port 4 nsew
flabel locali s 0 630 184 698 0 FreeSans 400 0 0 0 C2
port 5 nsew
flabel locali s 0 1070 184 1138 0 FreeSans 400 0 0 0 C4
port 6 nsew
flabel locali s 0 850 184 918 0 FreeSans 400 0 0 0 C8
port 7 nsew
flabel locali s 0 410 184 478 0 FreeSans 400 0 0 0 C16
port 8 nsew
<< end >>
