*RPLY_BIAS_SKY130A/RPLY_BIAS
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_BIAS_lpe.spi
#else
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_10_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_20_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHDLCM_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHL_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHDL_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_NCHDLCM_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_NCHDL_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_PCHDLA_lpe.spi
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_NCHL_lpe.spi
.include ../../../work/xsch/RPLY_BIAS.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter gmin=1e-12 method=gear
#else
.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter gmin=1e-15 method=gear
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param T_END = {10u}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc {AVDD}
VPWR  PWRUP_1V8  VSS  dc {AVDD}

*-----------------------------------------------------------------
* Middlebrook loop method
*-----------------------------------------------------------------
* V1 = Input to the feedback loop
* V2 = Output of the amplifier, or where you break the loop
* Middlebrook sources http://education.ingenazure.com/ac-stability-analysis-ngspice/
VLSTB1 LSTBPROBE LPI dc 0 ac 0
VLSTB2 LSTBPROBE LPO dc 0
ILSTB1 0 LSTBPROBE  dc 0 ac 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------

XDUT VDD_1V8 VSS PWRUP_1V8 LPI LPO
+ IBP_1U<3>,IBP_1U<2>,IBP_1U<1>,IBP_1U<0> T_OP T_ON RPLY_BIAS
*-----------------------------------------------------------------
* STASH
*-----------------------------------------------------------------

V3 IBP_1U<3> 0 dc {AVDD/2}
V2 IBP_1U<2> 0 dc {AVDD/2}
V1 IBP_1U<1> 0 dc {AVDD/2}
V0 IBP_1U<0> 0 dc {AVDD/2}


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save i(vlstb1) i(vlstb2) v(lstbprobe) v(LPO) v(LPI) v(xdut.vr1) v(xdut.vd1)
#ifdef Debug
*.save all
#else
*.probe v(VDD_1V8) v(VSS) v(PWRUP_1V8) v(LPI) v(LPO) v(IBP_1U) i(v1)
*+ v(XDUT.VD1) v(XDUT.VD2) v(XDUT.VR1) v(D_VD) v(D_VD_REF) v(D_VD_ERR)
*+ v(V_OFF) i(VDD)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
*pre_set strict_errorhandling
*pre_set ng_nomodcheck
set num_threads=8
set color0=white
set color1=black
unset askquit


optran 0 0 0 10n 1u 0

op
write {cicname}_op.raw


*----------------------------------------------------------------
* Middlebrook sources http://education.ingenazure.com/ac-stability-analysis-ngspice/
*----------------------------------------------------------------
* Set voltage AC to 1
alter @vlstb1[ac]=1
alter @ilstb1[ac]=0
ac dec 50 100 1T
write {cicname}_0.raw all

* Set Current to 1
alter @vlstb2[acmag]=0
alter @vlstb1[acmag]=1
ac dec 50 100 1T
write {cicname}_1.raw all




#ifdef Debug


*quit
#else

quit
#endif
.endc
