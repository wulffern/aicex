magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 2560
<< locali >>
rect 720 210 874 270
rect 720 370 874 430
rect 720 850 874 910
rect 720 1010 874 1070
rect 720 1490 874 1550
rect 720 1650 874 1710
rect 720 2130 874 2190
rect 720 2290 874 2350
rect 874 210 1380 270
rect 874 370 1380 430
rect 874 850 1380 910
rect 874 1010 1380 1070
rect 874 1490 1380 1550
rect 874 1650 1380 1710
rect 874 2130 1380 2190
rect 874 2290 1380 2350
rect 874 210 934 2350
rect 330 130 390 2430
rect 1710 130 1770 2430
rect 270 130 450 190
rect 630 210 810 270
rect 2010 120 2190 200
rect -90 120 90 200
<< poly >>
rect 270 142 1830 178
rect 270 462 1830 498
rect 270 782 1830 818
rect 270 1102 1830 1138
rect 270 1422 1830 1458
rect 270 1742 1830 1778
rect 270 2062 1830 2098
rect 270 2382 1830 2418
<< m3 >>
rect 1290 0 1474 2560
rect 630 0 814 2560
rect 1290 0 1474 2560
rect 630 0 814 2560
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1050 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1050 1280
use NCHDL MN4
transform 1 0 0 0 1 1280
box 0 1280 1050 1600
use NCHDL MN5
transform 1 0 0 0 1 1600
box 0 1600 1050 1920
use NCHDL MN6
transform 1 0 0 0 1 1920
box 0 1920 1050 2240
use NCHDL MN7
transform 1 0 0 0 1 2240
box 0 2240 1050 2560
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL MP2
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use PCHDL MP3
transform 1 0 1050 0 1 960
box 1050 960 2100 1280
use PCHDL MP4
transform 1 0 1050 0 1 1280
box 1050 1280 2100 1600
use PCHDL MP5
transform 1 0 1050 0 1 1600
box 1050 1600 2100 1920
use PCHDL MP6
transform 1 0 1050 0 1 1920
box 1050 1920 2100 2240
use PCHDL MP7
transform 1 0 1050 0 1 2240
box 1050 2240 2100 2560
use cut_M1M4_2x1 
transform 1 0 1290 0 1 50
box 1290 50 1474 118
use cut_M1M4_2x1 
transform 1 0 1290 0 1 530
box 1290 530 1474 598
use cut_M1M4_2x1 
transform 1 0 1290 0 1 690
box 1290 690 1474 758
use cut_M1M4_2x1 
transform 1 0 1290 0 1 1170
box 1290 1170 1474 1238
use cut_M1M4_2x1 
transform 1 0 1290 0 1 1330
box 1290 1330 1474 1398
use cut_M1M4_2x1 
transform 1 0 1290 0 1 1810
box 1290 1810 1474 1878
use cut_M1M4_2x1 
transform 1 0 1290 0 1 1970
box 1290 1970 1474 2038
use cut_M1M4_2x1 
transform 1 0 1290 0 1 2450
box 1290 2450 1474 2518
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M4_2x1 
transform 1 0 630 0 1 690
box 630 690 814 758
use cut_M1M4_2x1 
transform 1 0 630 0 1 1170
box 630 1170 814 1238
use cut_M1M4_2x1 
transform 1 0 630 0 1 1330
box 630 1330 814 1398
use cut_M1M4_2x1 
transform 1 0 630 0 1 1810
box 630 1810 814 1878
use cut_M1M4_2x1 
transform 1 0 630 0 1 1970
box 630 1970 814 2038
use cut_M1M4_2x1 
transform 1 0 630 0 1 2450
box 630 2450 814 2518
<< labels >>
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 630 210 810 270 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 3 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 4 nsew
flabel m3 s 1290 0 1474 2560 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 630 0 814 2560 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
