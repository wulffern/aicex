** sch_path:
*+ /Users/wulff/pro/aicex/ip/sun_pll_sky130nm/work/../design/SUN_PLL_SKY130NM/SUN_PLL_ROSC.sch
.subckt SUN_PLL_ROSC PWRUP_1V8 VDD_ROSC AVSS VDD_1V8 CK
*.ipin PWRUP_1V8
*.ipin VDD_ROSC
*.ipin AVSS
*.ipin VDD_1V8
*.opin CK
xa3 VDD_1V8 CKUP __UNCONNECTED_PIN__0 NI N_7 AVSS SUN_PLL_LSCORE
xa4 CKUP CK VDD_1V8 AVSS SUNTR_IVX1_CV
xa5 VDD_1V8 AVSS SUNTR_TAPCELLB_CV
xb1 PWRUP_1V8 N_0 NI VDD_ROSC AVSS SUNTR_NDX1_CV
xb2_0 N_1 N_0 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_1 N_2 N_1 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_2 N_3 N_2 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_3 N_4 N_3 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_4 N_5 N_4 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_5 N_6 N_5 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_6 N_7 N_6 VDD_ROSC AVSS SUNTR_IVX1_CV
xb2_7 NI N_7 VDD_ROSC AVSS SUNTR_IVX1_CV
.ends

* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sym # of pins=6
** sym_path:
*+ /Users/wulff/Documents/pro/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sym
** sch_path:
*+ /Users/wulff/Documents/pro/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sch
.subckt SUN_PLL_LSCORE  AVDD YN Y A AN AVSS
*.ipin AVDD
*.ipin A
*.ipin AN
*.opin Y
*.opin YN
*.ipin AVSS
xb1_0 Y AN AVSS AVSS SUNTR_NCHDL
xb1_1 Y AN AVSS AVSS SUNTR_NCHDL
xb2_0 YN A AVSS AVSS SUNTR_NCHDL
xb2_1 YN A AVSS AVSS SUNTR_NCHDL
xc1a net2 YN AVDD AVDD SUNTR_PCHDL
xc1b Y YN net2 AVDD SUNTR_PCHDL
xc2a net1 Y AVDD AVDD SUNTR_PCHDL
xc2b YN Y net1 AVDD SUNTR_PCHDL
.ends

.end
