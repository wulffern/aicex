magic
tech sky130A
magscale 1 2
timestamp 1658699483
<< checkpaint >>
rect -3928 -1848 28016 52422
<< m3 >>
rect 9100 28760 26178 28836
rect 9100 29148 26178 29224
rect 24104 29528 24180 37032
rect 24384 29528 24460 44776
rect 3944 29612 4020 40544
rect 4824 29806 4900 40544
rect 8984 30000 9060 40544
rect -216 30194 -140 40544
rect -216 30194 -140 40544
rect 13432 30388 13508 40570
rect 13432 30388 13508 40570
rect 18472 30582 18548 40570
rect 18472 30582 18548 40570
rect 10579 30776 10655 40570
rect 10579 30776 10655 40570
rect 15619 30970 15695 40570
rect 15619 30970 15695 40570
rect 499 31164 575 40570
rect 5539 31358 5615 40570
rect 5539 31358 5615 40570
rect 3352 31552 3428 40570
rect 3352 31552 3428 40570
rect 8392 31746 8468 40570
rect 8392 31746 8468 40570
rect 659 31940 735 41978
rect 8232 32134 8308 41978
rect 5699 32328 5775 41978
rect 3192 32522 3268 41978
rect 10914 32716 10990 43386
rect 13098 32910 13174 43386
rect 15954 33104 16030 43386
rect 8058 33298 8134 43386
rect 3018 33492 3094 43386
rect 834 33686 910 43386
rect 18138 33880 18214 43386
rect 5874 34074 5950 43386
rect 200 34774 400 50982
rect 3528 34774 3728 50982
rect 5240 34774 5440 50982
rect 8568 34774 8768 50982
rect 10280 34774 10480 50982
rect 13608 34774 13808 50982
rect 15320 34774 15520 50982
rect 18648 34774 18848 50982
rect 20360 34774 20560 50982
rect 23688 34774 23888 50982
rect 9648 -720 9848 5280
rect 14240 -720 14440 5280
rect 992 34774 1192 51702
rect 2736 34774 2936 51702
rect 6032 34774 6232 51702
rect 7776 34774 7976 51702
rect 11072 34774 11272 51702
rect 12816 34774 13016 51702
rect 16112 34774 16312 51702
rect 17856 34774 18056 51702
rect 21152 34774 21352 51702
rect 22896 34774 23096 51702
rect 8856 -1440 9056 5280
rect 15032 -1440 15232 5280
rect 1568 39584 1768 52422
rect 2160 39584 2360 52422
rect 6608 39584 6808 52422
rect 7200 39584 7400 52422
rect 11648 39584 11848 52422
rect 12240 39584 12440 52422
rect 16688 39584 16888 52422
rect 17280 39584 17480 52422
rect 21728 39584 21928 52422
rect 10294 -1848 10370 3470
rect 13718 -1848 13794 3470
rect 10924 1290 11180 1366
rect 9138 5474 10924 5550
rect 12908 1290 13088 1366
rect 13088 5474 14910 5550
rect 11180 1290 11360 1366
rect 11360 2698 12908 2774
rect 11360 1290 11436 2774
rect 11072 50 11272 126
rect 12816 50 13016 126
rect 20659 40570 20735 40770
<< m2 >>
rect 14872 28254 14948 28836
rect 9100 28254 9176 29224
rect 3944 29536 14020 29612
rect 4824 29730 13660 29806
rect 8984 29924 13300 30000
rect -216 30118 14380 30194
rect 11304 30312 13508 30388
rect 11664 30506 18548 30582
rect 10579 30700 11200 30776
rect 11484 30894 15695 30970
rect 499 31088 9760 31164
rect 5539 31282 10480 31358
rect 3352 31476 10120 31552
rect 8392 31670 10840 31746
rect 659 31864 9940 31940
rect 8232 32058 11020 32134
rect 5699 32252 10660 32328
rect 3192 32446 10300 32522
rect 10914 32640 12940 32716
rect 12684 32834 13174 32910
rect 12504 33028 16030 33104
rect 8058 33222 13120 33298
rect 3018 33416 13840 33492
rect 834 33610 14200 33686
rect 12324 33804 18214 33880
rect 5874 33998 13480 34074
rect 992 48766 1336 48842
rect 1336 48156 3944 48232
rect 3868 48156 3944 48356
rect 1336 48156 1412 48850
rect 6032 48766 6376 48842
rect 6376 48156 8984 48232
rect 8908 48156 8984 48356
rect 6376 48156 6452 48850
rect 11072 48766 11416 48842
rect 11416 48156 14024 48232
rect 13948 48156 14024 48356
rect 11416 48156 11492 48850
rect 16112 48766 16456 48842
rect 16456 48156 19064 48232
rect 18988 48156 19064 48356
rect 16456 48156 16532 48850
rect -232 44988 20144 45064
rect -308 44988 -232 45188
rect 3868 44988 3944 45188
rect 4732 44988 4808 45188
rect 8908 44988 8984 45188
rect 9772 44988 9848 45188
rect 13948 44988 14024 45188
rect 14812 44988 14888 45188
rect 18988 44988 19064 45188
rect 19852 44988 19928 45188
rect 1008 35528 1336 35604
rect 1336 35124 3944 35200
rect 3868 35124 3944 35340
rect 1336 35124 1412 35604
rect 6048 35528 6376 35604
rect 6376 35124 8984 35200
rect 8908 35124 8984 35340
rect 6376 35124 6452 35604
rect 11088 35528 11416 35604
rect 11416 35124 14024 35200
rect 13948 35124 14024 35340
rect 11416 35124 11492 35604
rect 16128 35528 16456 35604
rect 16456 35124 19064 35200
rect 18988 35124 19064 35340
rect 16456 35124 16532 35604
rect 21168 35528 21496 35604
rect 21496 35528 21572 35604
rect 2720 35528 3048 35604
rect 3048 35528 3124 35668
rect 3048 35668 4824 35744
rect 4748 35264 4824 35744
rect 7760 35528 8088 35604
rect 8088 35528 8164 35668
rect 8088 35668 9864 35744
rect 9788 35264 9864 35744
rect 12800 35528 13128 35604
rect 13128 35528 13204 35668
rect 13128 35668 14904 35744
rect 14828 35264 14904 35744
rect 17840 35528 18168 35604
rect 18168 35528 18244 35668
rect 18168 35668 19944 35744
rect 19868 35264 19944 35744
rect -216 37316 20144 37392
rect -292 37024 -216 37392
rect 3868 37024 3944 37392
rect 4748 37024 4824 37392
rect 8908 37024 8984 37392
rect 9788 37024 9864 37392
rect 13948 37024 14024 37392
rect 14828 37024 14904 37392
rect 18988 37024 19064 37392
rect 19868 37024 19944 37392
rect -232 37796 20144 37872
rect -308 37796 -232 38148
rect 3868 37796 3944 38148
rect 4732 37796 4808 38148
rect 8908 37796 8984 38148
rect 9772 37796 9848 38148
rect 13948 37796 14024 38148
rect 14812 37796 14888 38148
rect 18988 37796 19064 38148
rect 19852 37796 19928 38148
rect -16 38792 1424 38852
rect 1424 38792 1640 38852
rect 1424 38792 2504 38852
rect 1424 38792 6680 38852
rect 1424 38792 7544 38852
rect 1424 38792 11720 38852
rect 1424 38792 12584 38852
rect 1424 38792 16760 38852
rect 1424 38792 17624 38852
rect 1424 38792 21800 38852
rect 23396 40318 23780 40394
rect 20084 37100 23396 37176
rect 23396 37100 23472 40402
rect 20044 37024 20144 37100
rect 22740 41726 22988 41802
rect 20084 38164 22740 38240
rect 22740 38164 22816 41810
rect 20036 38088 20144 38164
rect 22556 49000 22728 49076
rect 20036 45832 22728 45908
rect 22728 45832 22804 49076
rect 22308 49704 22556 49780
rect 21260 48766 22308 48842
rect 22308 48766 22384 49780
rect 11180 2698 11352 2774
rect 11352 1290 12908 1366
rect 11352 1290 11428 2774
rect -232 38792 1640 38852
<< m4 >>
rect 24104 29148 24180 29528
rect 24384 28760 24460 29528
rect 10924 1290 11000 5550
rect 13088 1290 13164 5550
<< m1 >>
rect 13944 28194 14020 29536
rect 13584 28194 13660 29730
rect 13224 28194 13300 29924
rect 14304 28194 14380 30118
rect 11304 28194 11380 30312
rect 11664 28194 11740 30506
rect 11124 28194 11200 30700
rect 11484 28194 11560 30894
rect 9684 28194 9760 31088
rect 10404 28194 10480 31282
rect 10044 28194 10120 31476
rect 10764 28194 10840 31670
rect 9864 28194 9940 31864
rect 10944 28194 11020 32058
rect 10584 28194 10660 32252
rect 10224 28194 10300 32446
rect 12864 28194 12940 32640
rect 12684 28194 12760 32834
rect 12504 28194 12580 33028
rect 13044 28194 13120 33222
rect 13764 28194 13840 33416
rect 14124 28194 14200 33610
rect 12324 28194 12400 33804
rect 13404 28194 13480 33998
rect 10142 -1644 10202 558
rect 13886 -1644 13946 558
rect -3868 48296 -232 48356
rect 2720 48736 3056 48796
rect 3056 48176 4808 48236
rect 4748 48176 4808 48356
rect 3056 48176 3116 48804
rect 7760 48736 8096 48796
rect 8096 48176 9848 48236
rect 9788 48176 9848 48356
rect 8096 48176 8156 48804
rect 12800 48736 13136 48796
rect 13136 48176 14888 48236
rect 14828 48176 14888 48356
rect 13136 48176 13196 48804
rect 17840 48736 18176 48796
rect 18176 48176 19928 48236
rect 19868 48176 19928 48356
rect 18176 48176 18236 48804
rect 22328 49352 22556 49412
rect 20468 46624 22328 46684
rect 22328 46624 22388 49420
rect -3004 5474 76 5534
rect -3004 8314 76 8374
rect -3004 11154 76 11214
rect -3004 13994 76 14054
rect -3004 16834 76 16894
rect -3004 19674 76 19734
rect -3004 22514 76 22574
rect -3004 25354 76 25414
rect 23972 5474 27092 5534
rect 23972 8314 27092 8374
rect 23972 11154 27092 11214
rect 23972 13994 27092 14054
rect 23972 16834 27092 16894
rect 23972 19674 27092 19734
rect 23972 22514 27092 22574
rect 23972 25354 27092 25414
<< locali >>
rect 26892 -720 27092 50982
rect -3004 -720 27092 -520
rect -3004 50782 27092 50982
rect -3004 -720 -2804 50982
rect 26892 -720 27092 50982
rect 27612 -1440 27812 51702
rect -3724 -1440 27812 -1240
rect -3724 51502 27812 51702
rect -3724 -1440 -3524 51702
rect 27612 -1440 27812 51702
rect -3724 52222 27812 52422
rect -3724 52222 27812 52422
rect 27956 -1644 28016 52422
rect -3724 -1644 28016 -1584
rect 27956 -1644 28016 52422
rect -3928 -1848 28016 -1788
rect -3928 -1848 -3868 52422
rect 20360 46624 20576 46684
rect -232 45128 -16 45188
rect 1424 38792 1640 38852
rect 11072 2698 11288 2758
rect 11072 1290 11288 1350
use SARBSSW_CV XB1
transform -1 0 12044 0 1 0
box 12044 0 26372 5280
use SARBSSW_CV XB2
transform 1 0 12044 0 1 0
box 12044 0 26372 5280
use CDAC8_CV XDAC1
transform -1 0 11844 0 1 5474
box 11844 5474 23576 28254
use CDAC8_CV XDAC2
transform 1 0 12204 0 1 5474
box 12204 5474 23936 28254
use SARDIGEX4_CV XA0
transform 1 0 -556 0 1 34774
box -556 34774 1964 49206
use SARDIGEX4_CV XA1
transform -1 0 4484 0 1 34774
box 4484 34774 7004 49206
use SARDIGEX4_CV XA2
transform 1 0 4484 0 1 34774
box 4484 34774 7004 49206
use SARDIGEX4_CV XA3
transform -1 0 9524 0 1 34774
box 9524 34774 12044 49206
use SARDIGEX4_CV XA4
transform 1 0 9524 0 1 34774
box 9524 34774 12044 49206
use SARDIGEX4_CV XA5
transform -1 0 14564 0 1 34774
box 14564 34774 17084 49206
use SARDIGEX4_CV XA6
transform 1 0 14564 0 1 34774
box 14564 34774 17084 49206
use SARDIGEX4_CV XA7
transform -1 0 19604 0 1 34774
box 19604 34774 22124 49206
use SARDIGEX4_CV XA8
transform 1 0 19604 0 1 34774
box 19604 34774 22124 49206
use SARCMPX1_CV XA20
transform -1 0 24644 0 1 34774
box 24644 34774 27164 50262
use cut_M3M4_1x2 
transform 1 0 14872 0 1 28254
box 14872 28254 14948 28454
use cut_M3M4_2x1 
transform 1 0 14872 0 1 28760
box 14872 28760 15072 28836
use cut_M3M4_1x2 
transform 1 0 9100 0 1 28254
box 9100 28254 9176 28454
use cut_M3M4_2x1 
transform 1 0 9100 0 1 29148
box 9100 29148 9300 29224
use cut_M2M4_2x1 
transform 1 0 24104 0 1 37032
box 24104 37032 24304 37108
use cut_M4M5_2x1 
transform 1 0 24104 0 1 29148
box 24104 29148 24304 29224
use cut_M4M5_1x2 
transform 1 0 24104 0 1 29528
box 24104 29528 24180 29728
use cut_M3M4_2x1 
transform 1 0 24260 0 1 44776
box 24260 44776 24460 44852
use cut_M2M3_2x1 
transform 1 0 24104 0 1 44776
box 24104 44776 24304 44852
use cut_M4M5_2x1 
transform 1 0 24384 0 1 28760
box 24384 28760 24584 28836
use cut_M4M5_1x2 
transform 1 0 24384 0 1 29528
box 24384 29528 24460 29728
use cut_M3M4_1x2 
transform 1 0 3944 0 1 29474
box 3944 29474 4020 29674
use cut_M2M3_1x2 
transform 1 0 13936 0 1 29474
box 13936 29474 14012 29674
use cut_M3M4_1x2 
transform 1 0 4824 0 1 29668
box 4824 29668 4900 29868
use cut_M2M3_1x2 
transform 1 0 13576 0 1 29668
box 13576 29668 13652 29868
use cut_M3M4_1x2 
transform 1 0 8984 0 1 29862
box 8984 29862 9060 30062
use cut_M2M3_1x2 
transform 1 0 13216 0 1 29862
box 13216 29862 13292 30062
use cut_M3M4_1x2 
transform 1 0 -216 0 1 30056
box -216 30056 -140 30256
use cut_M2M3_1x2 
transform 1 0 14296 0 1 30056
box 14296 30056 14372 30256
use cut_M3M4_1x2 
transform 1 0 13432 0 1 30250
box 13432 30250 13508 30450
use cut_M2M3_1x2 
transform 1 0 11296 0 1 30250
box 11296 30250 11372 30450
use cut_M3M4_1x2 
transform 1 0 18472 0 1 30444
box 18472 30444 18548 30644
use cut_M2M3_1x2 
transform 1 0 11656 0 1 30444
box 11656 30444 11732 30644
use cut_M3M4_1x2 
transform 1 0 10579 0 1 30638
box 10579 30638 10655 30838
use cut_M2M3_1x2 
transform 1 0 11116 0 1 30638
box 11116 30638 11192 30838
use cut_M3M4_1x2 
transform 1 0 15619 0 1 30832
box 15619 30832 15695 31032
use cut_M2M3_1x2 
transform 1 0 11476 0 1 30832
box 11476 30832 11552 31032
use cut_M3M4_1x2 
transform 1 0 499 0 1 31026
box 499 31026 575 31226
use cut_M2M3_1x2 
transform 1 0 9676 0 1 31026
box 9676 31026 9752 31226
use cut_M3M4_1x2 
transform 1 0 5539 0 1 31220
box 5539 31220 5615 31420
use cut_M2M3_1x2 
transform 1 0 10396 0 1 31220
box 10396 31220 10472 31420
use cut_M3M4_1x2 
transform 1 0 3352 0 1 31414
box 3352 31414 3428 31614
use cut_M2M3_1x2 
transform 1 0 10036 0 1 31414
box 10036 31414 10112 31614
use cut_M3M4_1x2 
transform 1 0 8392 0 1 31608
box 8392 31608 8468 31808
use cut_M2M3_1x2 
transform 1 0 10756 0 1 31608
box 10756 31608 10832 31808
use cut_M3M4_1x2 
transform 1 0 659 0 1 31802
box 659 31802 735 32002
use cut_M2M3_1x2 
transform 1 0 9856 0 1 31802
box 9856 31802 9932 32002
use cut_M3M4_1x2 
transform 1 0 8232 0 1 31996
box 8232 31996 8308 32196
use cut_M2M3_1x2 
transform 1 0 10936 0 1 31996
box 10936 31996 11012 32196
use cut_M3M4_1x2 
transform 1 0 5699 0 1 32190
box 5699 32190 5775 32390
use cut_M2M3_1x2 
transform 1 0 10576 0 1 32190
box 10576 32190 10652 32390
use cut_M3M4_1x2 
transform 1 0 3192 0 1 32384
box 3192 32384 3268 32584
use cut_M2M3_1x2 
transform 1 0 10216 0 1 32384
box 10216 32384 10292 32584
use cut_M3M4_1x2 
transform 1 0 10914 0 1 32578
box 10914 32578 10990 32778
use cut_M2M3_1x2 
transform 1 0 12856 0 1 32578
box 12856 32578 12932 32778
use cut_M3M4_1x2 
transform 1 0 13098 0 1 32772
box 13098 32772 13174 32972
use cut_M2M3_1x2 
transform 1 0 12676 0 1 32772
box 12676 32772 12752 32972
use cut_M3M4_1x2 
transform 1 0 15954 0 1 32966
box 15954 32966 16030 33166
use cut_M2M3_1x2 
transform 1 0 12496 0 1 32966
box 12496 32966 12572 33166
use cut_M3M4_1x2 
transform 1 0 8058 0 1 33160
box 8058 33160 8134 33360
use cut_M2M3_1x2 
transform 1 0 13036 0 1 33160
box 13036 33160 13112 33360
use cut_M3M4_1x2 
transform 1 0 3018 0 1 33354
box 3018 33354 3094 33554
use cut_M2M3_1x2 
transform 1 0 13756 0 1 33354
box 13756 33354 13832 33554
use cut_M3M4_1x2 
transform 1 0 834 0 1 33548
box 834 33548 910 33748
use cut_M2M3_1x2 
transform 1 0 14116 0 1 33548
box 14116 33548 14192 33748
use cut_M3M4_1x2 
transform 1 0 18138 0 1 33742
box 18138 33742 18214 33942
use cut_M2M3_1x2 
transform 1 0 12316 0 1 33742
box 12316 33742 12392 33942
use cut_M3M4_1x2 
transform 1 0 5874 0 1 33936
box 5874 33936 5950 34136
use cut_M2M3_1x2 
transform 1 0 13396 0 1 33936
box 13396 33936 13472 34136
use cut_M1M4_2x2 
transform 1 0 200 0 1 50782
box 200 50782 400 50982
use cut_M1M4_2x2 
transform 1 0 3528 0 1 50782
box 3528 50782 3728 50982
use cut_M1M4_2x2 
transform 1 0 5240 0 1 50782
box 5240 50782 5440 50982
use cut_M1M4_2x2 
transform 1 0 8568 0 1 50782
box 8568 50782 8768 50982
use cut_M1M4_2x2 
transform 1 0 10280 0 1 50782
box 10280 50782 10480 50982
use cut_M1M4_2x2 
transform 1 0 13608 0 1 50782
box 13608 50782 13808 50982
use cut_M1M4_2x2 
transform 1 0 15320 0 1 50782
box 15320 50782 15520 50982
use cut_M1M4_2x2 
transform 1 0 18648 0 1 50782
box 18648 50782 18848 50982
use cut_M1M4_2x2 
transform 1 0 20360 0 1 50782
box 20360 50782 20560 50982
use cut_M1M4_2x2 
transform 1 0 23688 0 1 50782
box 23688 50782 23888 50982
use cut_M1M4_2x2 
transform 1 0 9648 0 1 -720
box 9648 -720 9848 -520
use cut_M1M4_2x2 
transform 1 0 14240 0 1 -720
box 14240 -720 14440 -520
use cut_M1M4_2x2 
transform 1 0 992 0 1 51502
box 992 51502 1192 51702
use cut_M1M4_2x2 
transform 1 0 2736 0 1 51502
box 2736 51502 2936 51702
use cut_M1M4_2x2 
transform 1 0 6032 0 1 51502
box 6032 51502 6232 51702
use cut_M1M4_2x2 
transform 1 0 7776 0 1 51502
box 7776 51502 7976 51702
use cut_M1M4_2x2 
transform 1 0 11072 0 1 51502
box 11072 51502 11272 51702
use cut_M1M4_2x2 
transform 1 0 12816 0 1 51502
box 12816 51502 13016 51702
use cut_M1M4_2x2 
transform 1 0 16112 0 1 51502
box 16112 51502 16312 51702
use cut_M1M4_2x2 
transform 1 0 17856 0 1 51502
box 17856 51502 18056 51702
use cut_M1M4_2x2 
transform 1 0 21152 0 1 51502
box 21152 51502 21352 51702
use cut_M1M4_2x2 
transform 1 0 22896 0 1 51502
box 22896 51502 23096 51702
use cut_M1M4_2x2 
transform 1 0 8856 0 1 -1440
box 8856 -1440 9056 -1240
use cut_M1M4_2x2 
transform 1 0 15032 0 1 -1440
box 15032 -1440 15232 -1240
use cut_M1M4_2x2 
transform 1 0 1568 0 1 52222
box 1568 52222 1768 52422
use cut_M1M4_2x2 
transform 1 0 2160 0 1 52222
box 2160 52222 2360 52422
use cut_M1M4_2x2 
transform 1 0 6608 0 1 52222
box 6608 52222 6808 52422
use cut_M1M4_2x2 
transform 1 0 7200 0 1 52222
box 7200 52222 7400 52422
use cut_M1M4_2x2 
transform 1 0 11648 0 1 52222
box 11648 52222 11848 52422
use cut_M1M4_2x2 
transform 1 0 12240 0 1 52222
box 12240 52222 12440 52422
use cut_M1M4_2x2 
transform 1 0 16688 0 1 52222
box 16688 52222 16888 52422
use cut_M1M4_2x2 
transform 1 0 17280 0 1 52222
box 17280 52222 17480 52422
use cut_M1M4_2x2 
transform 1 0 21728 0 1 52222
box 21728 52222 21928 52422
use cut_M1M2_2x1 
transform 1 0 10080 0 1 498
box 10080 498 10264 566
use cut_M1M2_2x1 
transform 1 0 10080 0 1 -1644
box 10080 -1644 10264 -1576
use cut_M1M2_2x1 
transform 1 0 13824 0 1 498
box 13824 498 14008 566
use cut_M1M2_2x1 
transform 1 0 13824 0 1 -1644
box 13824 -1644 14008 -1576
use cut_M1M2_2x1 
transform 1 0 -232 0 1 48296
box -232 48296 -48 48364
use cut_M1M2_1x2 
transform 1 0 -3932 0 1 48234
box -3932 48234 -3864 48418
use cut_M1M4_2x1 
transform 1 0 10232 0 1 -1848
box 10232 -1848 10432 -1772
use cut_M1M4_2x1 
transform 1 0 13656 0 1 -1848
box 13656 -1848 13856 -1772
use cut_M1M3_2x1 
transform 1 0 992 0 1 48774
box 992 48774 1192 48850
use cut_M1M3_2x1 
transform 1 0 3944 0 1 48296
box 3944 48296 4144 48372
use cut_M1M3_2x1 
transform 1 0 6032 0 1 48774
box 6032 48774 6232 48850
use cut_M1M3_2x1 
transform 1 0 8984 0 1 48296
box 8984 48296 9184 48372
use cut_M1M3_2x1 
transform 1 0 11072 0 1 48774
box 11072 48774 11272 48850
use cut_M1M3_2x1 
transform 1 0 14024 0 1 48296
box 14024 48296 14224 48372
use cut_M1M3_2x1 
transform 1 0 16112 0 1 48774
box 16112 48774 16312 48850
use cut_M1M3_2x1 
transform 1 0 19064 0 1 48296
box 19064 48296 19264 48372
use cut_M1M3_2x1 
transform 1 0 -232 0 1 45128
box -232 45128 -32 45204
use cut_M1M3_2x1 
transform 1 0 3944 0 1 45128
box 3944 45128 4144 45204
use cut_M1M3_2x1 
transform 1 0 4808 0 1 45128
box 4808 45128 5008 45204
use cut_M1M3_2x1 
transform 1 0 8984 0 1 45128
box 8984 45128 9184 45204
use cut_M1M3_2x1 
transform 1 0 9848 0 1 45128
box 9848 45128 10048 45204
use cut_M1M3_2x1 
transform 1 0 14024 0 1 45128
box 14024 45128 14224 45204
use cut_M1M3_2x1 
transform 1 0 14888 0 1 45128
box 14888 45128 15088 45204
use cut_M1M3_2x1 
transform 1 0 19064 0 1 45128
box 19064 45128 19264 45204
use cut_M1M3_2x1 
transform 1 0 19928 0 1 45128
box 19928 45128 20128 45204
use cut_M1M2_2x1 
transform 1 0 2720 0 1 48736
box 2720 48736 2904 48804
use cut_M1M2_2x1 
transform 1 0 4808 0 1 48296
box 4808 48296 4992 48364
use cut_M1M2_2x1 
transform 1 0 7760 0 1 48736
box 7760 48736 7944 48804
use cut_M1M2_2x1 
transform 1 0 9848 0 1 48296
box 9848 48296 10032 48364
use cut_M1M2_2x1 
transform 1 0 12800 0 1 48736
box 12800 48736 12984 48804
use cut_M1M2_2x1 
transform 1 0 14888 0 1 48296
box 14888 48296 15072 48364
use cut_M1M2_2x1 
transform 1 0 17840 0 1 48736
box 17840 48736 18024 48804
use cut_M1M2_2x1 
transform 1 0 19928 0 1 48296
box 19928 48296 20112 48364
use cut_M1M3_2x1 
transform 1 0 -232 0 1 38088
box -232 38088 -32 38164
use cut_M1M3_2x1 
transform 1 0 3944 0 1 38088
box 3944 38088 4144 38164
use cut_M1M3_2x1 
transform 1 0 4808 0 1 38088
box 4808 38088 5008 38164
use cut_M1M3_2x1 
transform 1 0 8984 0 1 38088
box 8984 38088 9184 38164
use cut_M1M3_2x1 
transform 1 0 9848 0 1 38088
box 9848 38088 10048 38164
use cut_M1M3_2x1 
transform 1 0 14024 0 1 38088
box 14024 38088 14224 38164
use cut_M1M3_2x1 
transform 1 0 14888 0 1 38088
box 14888 38088 15088 38164
use cut_M1M3_2x1 
transform 1 0 19064 0 1 38088
box 19064 38088 19264 38164
use cut_M1M3_2x1 
transform 1 0 19928 0 1 38088
box 19928 38088 20128 38164
use cut_M1M3_2x1 
transform 1 0 1424 0 1 38792
box 1424 38792 1624 38868
use cut_M1M3_2x1 
transform 1 0 1424 0 1 38792
box 1424 38792 1624 38868
use cut_M1M3_2x1 
transform 1 0 2288 0 1 38792
box 2288 38792 2488 38868
use cut_M1M3_2x1 
transform 1 0 6464 0 1 38792
box 6464 38792 6664 38868
use cut_M1M3_2x1 
transform 1 0 7328 0 1 38792
box 7328 38792 7528 38868
use cut_M1M3_2x1 
transform 1 0 11504 0 1 38792
box 11504 38792 11704 38868
use cut_M1M3_2x1 
transform 1 0 12368 0 1 38792
box 12368 38792 12568 38868
use cut_M1M3_2x1 
transform 1 0 16544 0 1 38792
box 16544 38792 16744 38868
use cut_M1M3_2x1 
transform 1 0 17408 0 1 38792
box 17408 38792 17608 38868
use cut_M1M3_2x1 
transform 1 0 21584 0 1 38792
box 21584 38792 21784 38868
use cut_M1M3_2x1 
transform 1 0 23688 0 1 40326
box 23688 40326 23888 40402
use cut_M1M3_2x1 
transform 1 0 22896 0 1 41734
box 22896 41734 23096 41810
use cut_M1M3_2x1 
transform 1 0 22448 0 1 49000
box 22448 49000 22648 49076
use cut_M1M3_2x1 
transform 1 0 19928 0 1 45832
box 19928 45832 20128 45908
use cut_M1M3_2x1 
transform 1 0 22464 0 1 49704
box 22464 49704 22664 49780
use cut_M1M3_2x1 
transform 1 0 21168 0 1 48774
box 21168 48774 21368 48850
use cut_M1M2_2x1 
transform 1 0 22480 0 1 49352
box 22480 49352 22664 49420
use cut_M1M2_2x1 
transform 1 0 20392 0 1 46624
box 20392 46624 20576 46692
use cut_M4M5_1x2 
transform 1 0 10924 0 1 1290
box 10924 1290 11000 1490
use cut_M4M5_1x2 
transform 1 0 10924 0 1 5350
box 10924 5350 11000 5550
use cut_M1M4_2x1 
transform 1 0 12800 0 1 1290
box 12800 1290 13000 1366
use cut_M4M5_1x2 
transform 1 0 13088 0 1 1290
box 13088 1290 13164 1490
use cut_M4M5_1x2 
transform 1 0 13088 0 1 5350
box 13088 5350 13164 5550
use cut_M1M3_2x1 
transform 1 0 11072 0 1 2698
box 11072 2698 11272 2774
use cut_M1M3_2x1 
transform 1 0 12800 0 1 1290
box 12800 1290 13000 1366
use cut_M1M4_2x1 
transform 1 0 11072 0 1 1290
box 11072 1290 11272 1366
use cut_M1M4_2x1 
transform 1 0 12800 0 1 2698
box 12800 2698 13000 2774
use cut_M1M3_2x1 
transform 1 0 -232 0 1 38792
box -232 38792 -32 38868
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 5534
box -3004 5534 -2820 5718
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 8374
box -3004 8374 -2820 8558
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 11214
box -3004 11214 -2820 11398
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 14054
box -3004 14054 -2820 14238
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 16894
box -3004 16894 -2820 17078
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 19734
box -3004 19734 -2820 19918
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 22574
box -3004 22574 -2820 22758
use cut_M1M2_2x2 
transform 1 0 -3004 0 1 25414
box -3004 25414 -2820 25598
use cut_M1M2_2x2 
transform 1 0 26908 0 1 5474
box 26908 5474 27092 5658
use cut_M1M2_2x2 
transform 1 0 26908 0 1 8314
box 26908 8314 27092 8498
use cut_M1M2_2x2 
transform 1 0 26908 0 1 11154
box 26908 11154 27092 11338
use cut_M1M2_2x2 
transform 1 0 26908 0 1 13994
box 26908 13994 27092 14178
use cut_M1M2_2x2 
transform 1 0 26908 0 1 16834
box 26908 16834 27092 17018
use cut_M1M2_2x2 
transform 1 0 26908 0 1 19674
box 26908 19674 27092 19858
use cut_M1M2_2x2 
transform 1 0 26908 0 1 22514
box 26908 22514 27092 22698
use cut_M1M2_2x2 
transform 1 0 26908 0 1 25354
box 26908 25354 27092 25538
<< labels >>
flabel m3 s -216 30194 -140 40544 0 FreeSans 400 0 0 0 D<8>
port 6 nsew
flabel m3 s 13432 30388 13508 40570 0 FreeSans 400 0 0 0 D<3>
port 11 nsew
flabel m3 s 18472 30582 18548 40570 0 FreeSans 400 0 0 0 D<1>
port 13 nsew
flabel m3 s 10579 30776 10655 40570 0 FreeSans 400 0 0 0 D<4>
port 10 nsew
flabel m3 s 15619 30970 15695 40570 0 FreeSans 400 0 0 0 D<2>
port 12 nsew
flabel m3 s 5539 31358 5615 40570 0 FreeSans 400 0 0 0 D<6>
port 8 nsew
flabel m3 s 3352 31552 3428 40570 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8392 31746 8468 40570 0 FreeSans 400 0 0 0 D<5>
port 9 nsew
flabel locali s 26892 -720 27092 50982 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
flabel locali s 27612 -1440 27812 51702 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel locali s -3724 52222 27812 52422 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel locali s 27956 -1644 28016 52422 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel locali s 20360 46624 20576 46684 0 FreeSans 400 0 0 0 DONE
port 5 nsew
flabel m3 s 11072 50 11272 126 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew
flabel m3 s 12816 50 13016 126 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew
flabel locali s -232 45128 -16 45188 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 1424 38792 1640 38852 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s 11072 2698 11288 2758 0 FreeSans 400 0 0 0 SARN
port 3 nsew
flabel locali s 11072 1290 11288 1350 0 FreeSans 400 0 0 0 SARP
port 4 nsew
flabel m3 s 20659 40570 20735 40770 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
<< end >>
