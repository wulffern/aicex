magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 4480
<< locali >>
rect 1260 210 1398 270
rect 1398 710 1590 770
rect 1398 210 1458 770
rect 1530 770 1620 830
rect 1260 850 1398 910
rect 1398 1410 1620 1470
rect 1398 3970 1620 4030
rect 1398 850 1458 4030
rect 360 2050 498 2110
rect 498 850 720 910
rect 498 850 558 2110
rect 390 2950 498 3010
rect 498 850 720 910
rect 498 850 558 3010
rect 360 3010 450 3070
rect 720 1490 858 1550
rect 720 2130 858 2190
rect 858 1490 918 2190
rect 360 4290 498 4350
rect 498 4050 720 4110
rect 498 4050 558 4350
<< m1 >>
rect 1620 2050 1758 2110
rect 1620 3010 1758 3070
rect 1260 210 1758 270
rect 1758 210 1818 3078
rect 390 1350 498 1410
rect 498 530 720 590
rect 498 530 558 1478
rect 360 1410 450 1470
rect 720 3090 858 3150
rect 720 4050 858 4110
rect 858 3090 918 4118
rect 360 2370 498 2430
rect 498 2130 720 2190
rect 498 2130 558 2438
rect 1260 2450 1398 2510
rect 1398 1730 1620 1790
rect 1398 2690 1620 2750
rect 1398 1730 1458 2758
rect 1260 4370 1398 4430
rect 1398 3650 1620 3710
rect 1398 3650 1458 4438
rect 162 450 360 510
rect 162 3330 360 3390
rect 162 450 222 3398
<< m2 >>
rect 360 3970 498 4030
rect 498 3010 1620 3070
rect 498 3010 558 4038
<< m3 >>
rect 1170 0 1354 4480
rect 630 0 814 4480
use NDX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 1980 640
use IVX1_CV XA2
transform 1 0 0 0 1 640
box 0 640 1980 960
use IVTRIX1_CV XA3
transform 1 0 0 0 1 960
box 0 960 1980 1600
use IVTRIX1_CV XA4
transform 1 0 0 0 1 1600
box 0 1600 1980 2240
use IVX1_CV XA5
transform 1 0 0 0 1 2240
box 0 2240 1980 2560
use IVTRIX1_CV XA6
transform 1 0 0 0 1 2560
box 0 2560 1980 3200
use NDTRIX1_CV XA7
transform 1 0 0 0 1 3200
box 0 3200 1980 4160
use IVX1_CV XA8
transform 1 0 0 0 1 4160
box 0 4160 1980 4480
use cut_M1M2_2x1 
transform 1 0 1530 0 1 2050
box 1530 2050 1714 2118
use cut_M1M2_2x1 
transform 1 0 1530 0 1 3010
box 1530 3010 1714 3078
use cut_M1M2_2x1 
transform 1 0 1170 0 1 210
box 1170 210 1354 278
use cut_M1M2_2x1 
transform 1 0 270 0 1 1410
box 270 1410 454 1478
use cut_M1M2_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M3_2x1 
transform 1 0 270 0 1 3970
box 270 3970 454 4038
use cut_M1M3_2x1 
transform 1 0 1530 0 1 3010
box 1530 3010 1714 3078
use cut_M1M2_2x1 
transform 1 0 630 0 1 3090
box 630 3090 814 3158
use cut_M1M2_2x1 
transform 1 0 630 0 1 4050
box 630 4050 814 4118
use cut_M1M2_2x1 
transform 1 0 270 0 1 2370
box 270 2370 454 2438
use cut_M1M2_2x1 
transform 1 0 630 0 1 2130
box 630 2130 814 2198
use cut_M1M2_2x1 
transform 1 0 1170 0 1 2450
box 1170 2450 1354 2518
use cut_M1M2_2x1 
transform 1 0 1530 0 1 1730
box 1530 1730 1714 1798
use cut_M1M2_2x1 
transform 1 0 1530 0 1 2690
box 1530 2690 1714 2758
use cut_M1M2_2x1 
transform 1 0 1170 0 1 4370
box 1170 4370 1354 4438
use cut_M1M2_2x1 
transform 1 0 1530 0 1 3650
box 1530 3650 1714 3718
use cut_M1M2_2x1 
transform 1 0 270 0 1 450
box 270 450 454 518
use cut_M1M2_2x1 
transform 1 0 270 0 1 3330
box 270 3330 454 3398
<< labels >>
flabel locali s 270 1090 450 1150 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 CK
port 2 nsew
flabel locali s 630 4370 810 4430 0 FreeSans 400 0 0 0 Q
port 3 nsew
flabel locali s 630 4050 810 4110 0 FreeSans 400 0 0 0 QN
port 4 nsew
flabel locali s 270 3330 450 3390 0 FreeSans 400 0 0 0 RN
port 5 nsew
flabel locali s 1890 120 2070 200 0 FreeSans 400 0 0 0 BULKP
port 6 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 7 nsew
flabel m3 s 1170 0 1354 4480 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 4480 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
