magic
tech sky130A
magscale 1 2
timestamp 1658775803
<< checkpaint >>
rect 0 0 2520 14432
<< locali >>
rect 432 5778 600 5838
rect 600 4458 864 4518
rect 600 4458 660 5838
rect 432 8594 600 8654
rect 600 7274 864 7334
rect 600 7274 660 8654
rect 1860 4370 2088 4430
rect 1656 4106 1860 4166
rect 1860 4106 1920 4430
rect 432 11762 600 11822
rect 600 11498 864 11558
rect 600 11498 660 11822
rect 402 11762 462 12174
rect 480 12758 600 12818
rect 600 12554 864 12614
rect 600 12554 660 12818
rect 480 12818 540 12878
rect 480 13110 600 13170
rect 600 12906 864 12966
rect 600 12906 660 13170
rect 480 13170 540 13230
rect 432 13874 600 13934
rect 600 13434 864 13494
rect 600 13434 660 13934
rect 1656 8682 1824 8742
rect 1824 10002 2088 10062
rect 1824 8682 1884 10062
rect 1980 4018 2196 4078
rect 324 3314 540 3374
rect 324 13522 540 13582
rect 1548 13962 1764 14022
rect 324 10354 540 10414
rect 756 11850 972 11910
<< m1 >>
rect 432 7186 600 7246
rect 600 3050 864 3110
rect 600 3050 660 7254
rect 2088 11410 2256 11470
rect 1656 762 2256 822
rect 2256 762 2316 11478
rect 432 12466 600 12526
rect 600 11146 864 11206
rect 600 11146 660 12534
rect 1656 5866 1824 5926
rect 1824 10706 2088 10766
rect 1824 5866 1884 10774
<< m3 >>
rect 2186 4810 2262 9234
rect 340 5770 540 5846
rect 1055 5796 1131 5996
rect 1215 7204 1291 7404
rect 1390 8612 1466 8812
rect 2124 4810 2324 5010
rect 1548 0 1748 14432
rect 756 0 956 14432
rect 1548 0 1748 14432
rect 756 0 956 14432
<< m2 >>
rect 340 2250 540 2326
rect 340 490 540 566
rect 1564 754 1764 830
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use SARMRYX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2520 4224
use SWX4_CV XA2
transform 1 0 0 0 1 4224
box 0 4224 2520 5632
use SWX4_CV XA3
transform 1 0 0 0 1 5632
box 0 5632 2520 7040
use SWX4_CV XA4
transform 1 0 0 0 1 7040
box 0 7040 2520 8448
use SWX4_CV XA5
transform 1 0 0 0 1 8448
box 0 8448 2520 9856
use SARCEX1_CV XA6
transform 1 0 0 0 1 9856
box 0 9856 2520 11264
use IVX1_CV XA7
transform 1 0 0 0 1 11264
box 0 11264 2520 11616
use IVX1_CV XA8
transform 1 0 0 0 1 11616
box 0 11616 2520 11968
use NDX1_CV XA9
transform 1 0 0 0 1 11968
box 0 11968 2520 12672
use IVX1_CV XA10
transform 1 0 0 0 1 12672
box 0 12672 2520 13024
use NRX1_CV XA11
transform 1 0 0 0 1 13024
box 0 13024 2520 13728
use IVX1_CV XA12
transform 1 0 0 0 1 13728
box 0 13728 2520 14080
use TAPCELLB_CV XA13
transform 1 0 0 0 1 14080
box 0 14080 2520 14432
use DMY_CV XA14
transform 1 0 0 0 1 14432
box 0 14432 0 14432
use cut_M1M2_2x1 
transform 1 0 324 0 1 7186
box 324 7186 508 7254
use cut_M1M2_2x1 
transform 1 0 756 0 1 3050
box 756 3050 940 3118
use cut_M1M2_2x1 
transform 1 0 1980 0 1 11410
box 1980 11410 2164 11478
use cut_M1M2_2x1 
transform 1 0 1548 0 1 762
box 1548 762 1732 830
use cut_M1M2_2x1 
transform 1 0 324 0 1 12466
box 324 12466 508 12534
use cut_M1M2_2x1 
transform 1 0 756 0 1 11146
box 756 11146 940 11214
use cut_M1M2_2x1 
transform 1 0 1548 0 1 5866
box 1548 5866 1732 5934
use cut_M1M2_2x1 
transform 1 0 1980 0 1 10706
box 1980 10706 2164 10774
use cut_M1M4_2x1 
transform 1 0 340 0 1 5770
box 340 5770 540 5846
use cut_M1M4_1x2 
transform 1 0 1055 0 1 5796
box 1055 5796 1131 5996
use cut_M1M4_1x2 
transform 1 0 1215 0 1 7204
box 1215 7204 1291 7404
use cut_M1M4_1x2 
transform 1 0 1390 0 1 8612
box 1390 8612 1466 8812
use cut_M2M3_2x1 
transform 1 0 1564 0 1 754
box 1564 754 1764 830
use cut_M2M3_2x1 
transform 1 0 340 0 1 490
box 340 490 540 566
use cut_M2M3_2x1 
transform 1 0 340 0 1 490
box 340 490 540 566
use cut_M2M3_2x1 
transform 1 0 340 0 1 2250
box 340 2250 540 2326
use cut_M2M3_2x1 
transform 1 0 340 0 1 2250
box 340 2250 540 2326
<< labels >>
flabel m2 s 340 2250 540 2326 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1980 4018 2196 4078 0 FreeSans 400 0 0 0 RST_N
port 4 nsew
flabel m2 s 340 490 540 566 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 324 3314 540 3374 0 FreeSans 400 0 0 0 CMP_ON
port 2 nsew
flabel m2 s 1564 754 1764 830 0 FreeSans 400 0 0 0 ENO
port 5 nsew
flabel m3 s 340 5770 540 5846 0 FreeSans 400 0 0 0 CN1
port 10 nsew
flabel m3 s 1055 5796 1131 5996 0 FreeSans 400 0 0 0 CP1
port 8 nsew
flabel m3 s 1215 7204 1291 7404 0 FreeSans 400 0 0 0 CP0
port 7 nsew
flabel m3 s 1390 8612 1466 8812 0 FreeSans 400 0 0 0 CN0
port 9 nsew
flabel locali s 324 13522 540 13582 0 FreeSans 400 0 0 0 CEIN
port 11 nsew
flabel locali s 1548 13962 1764 14022 0 FreeSans 400 0 0 0 CEO
port 12 nsew
flabel locali s 324 10354 540 10414 0 FreeSans 400 0 0 0 CKS
port 13 nsew
flabel locali s 756 11850 972 11910 0 FreeSans 400 0 0 0 DONE
port 6 nsew
flabel m3 s 2124 4810 2324 5010 0 FreeSans 400 0 0 0 VREF
port 14 nsew
flabel m3 s 1548 0 1748 14432 0 FreeSans 400 0 0 0 AVDD
port 15 nsew
flabel m3 s 756 0 956 14432 0 FreeSans 400 0 0 0 AVSS
port 16 nsew
<< end >>
