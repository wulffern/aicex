magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 43972 62648
<< locali >>
rect 43204 528 43444 62120
rect 528 528 43444 768
rect 528 61880 43444 62120
rect 528 528 768 62120
rect 43204 528 43444 62120
rect 43732 0 43972 62648
rect 0 0 43972 240
rect 0 62408 43972 62648
rect 0 0 240 62648
rect 43732 0 43972 62648
use SUN_PLL_PFD xaa0
transform 1 0 1056 0 1 1056
box 1056 1056 5112 6816
use SUN_PLL_CP xaa1
transform 1 0 5112 0 1 1056
box 5112 1056 9528 11744
use SUN_PLL_KICK xaa3
transform 1 0 9528 0 1 1056
box 9528 1056 13656 11568
use SUN_PLL_BUF xaa4
transform 1 0 13656 0 1 1056
box 13656 1056 18072 8752
use SUN_PLL_ROSC xaa5
transform 1 0 18072 0 1 1056
box 18072 1056 24648 6464
use SUN_PLL_DIVN xaa6
transform 1 0 24648 0 1 1056
box 24648 1056 38784 8092
use SUN_PLL_LPF xbb0
transform 1 0 1056 0 1 11744
box 1056 11744 40888 61592
use SUN_PLL_BIAS xbb1
transform 1 0 40888 0 1 11744
box 40888 11744 42916 30464
<< labels >>
flabel locali s 43204 528 43444 62120 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 43732 0 43972 62648 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
<< end >>
