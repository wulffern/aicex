magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 37816 26400
<< locali >>
rect 37576 0 37816 26400
rect 0 0 37816 240
rect 0 26160 37816 26400
rect 0 0 240 26400
rect 37576 0 37816 26400
rect 2986 21070 3310 21290
rect 826 3806 1150 4026
<< m3 >>
rect 20588 0 20804 280
rect 20696 200 37528 276
rect 20696 1160 37528 1236
rect 20696 2120 37528 2196
rect 20696 3080 37528 3156
rect 20696 4040 37528 4116
rect 20696 5000 37528 5076
rect 20696 5960 37528 6036
rect 20696 6920 37528 6996
rect 20696 7880 37528 7956
rect 20696 8840 37528 8916
rect 20696 9800 37528 9876
rect 20696 10760 37528 10836
rect 20696 11720 37528 11796
rect 20696 12680 37528 12756
rect 20696 13640 37528 13716
rect 20696 14600 37528 14676
rect 20696 15560 37528 15636
rect 20696 16520 37528 16596
rect 20696 17480 37528 17556
rect 20696 18440 37528 18516
rect 20696 19400 37528 19476
rect 20696 20360 37528 20436
rect 20696 21320 37528 21396
rect 20696 22280 37528 22356
rect 20696 23240 37528 23316
rect 20696 24200 37528 24276
rect 20696 25160 37528 25236
rect 37528 200 37604 25236
<< m1 >>
rect 988 8122 1270 8182
rect 1270 3806 3148 3866
rect 1270 3806 1330 8190
rect 988 16754 1414 16814
rect 1414 12438 3148 12498
rect 1414 12438 1474 16822
rect 3148 21070 3370 21130
rect 3370 3880 4036 3940
rect 3370 4840 4036 4900
rect 3370 5800 4036 5860
rect 3370 6760 4036 6820
rect 3370 7720 4036 7780
rect 3370 8680 4036 8740
rect 3370 9640 4036 9700
rect 3370 10600 4036 10660
rect 3370 11560 4036 11620
rect 3370 12520 4036 12580
rect 3370 13480 4036 13540
rect 3370 14440 4036 14500
rect 3370 15400 4036 15460
rect 3370 16360 4036 16420
rect 3370 17320 4036 17380
rect 3370 18280 4036 18340
rect 3370 19240 4036 19300
rect 3370 20200 4036 20260
rect 3370 21160 4036 21220
rect 3370 22120 4036 22180
rect 3370 23080 4036 23140
rect 3370 24040 4036 24100
rect 3370 25000 4036 25060
rect 3370 25960 4036 26020
rect 3370 3880 3430 26036
<< m2 >>
rect 988 12438 1278 12514
rect 1278 8122 3148 8198
rect 1278 8122 1354 12514
rect 988 21070 1566 21146
rect 1566 16754 3148 16830
rect 1566 16754 1642 21146
rect 988 3806 1214 3882
rect 1214 1000 4036 1076
rect 1214 1960 4036 2036
rect 1214 2920 4036 2996
rect 1214 1000 1290 3882
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa10
transform 1 0 240 0 1 416
box 240 416 3896 4556
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa20
transform 1 0 240 0 1 4732
box 240 4732 3896 8872
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa30
transform 1 0 240 0 1 9048
box 240 9048 3896 13188
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa40
transform 1 0 240 0 1 13364
box 240 13364 3896 17504
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa50
transform 1 0 240 0 1 17680
box 240 17680 3896 21820
use CAP_LPF xb10
transform -1 0 37576 0 1 240
box 37576 240 71256 1200
use CAP_LPF xb20
transform -1 0 37576 0 1 1200
box 37576 1200 71256 2160
use CAP_LPF xb21
transform -1 0 37576 0 1 2160
box 37576 2160 71256 3120
use CAP_LPF xb30
transform -1 0 37576 0 1 3120
box 37576 3120 71256 4080
use CAP_LPF xb31
transform -1 0 37576 0 1 4080
box 37576 4080 71256 5040
use CAP_LPF xb32
transform -1 0 37576 0 1 5040
box 37576 5040 71256 6000
use CAP_LPF xb33
transform -1 0 37576 0 1 6000
box 37576 6000 71256 6960
use CAP_LPF xb34
transform -1 0 37576 0 1 6960
box 37576 6960 71256 7920
use CAP_LPF xb35
transform -1 0 37576 0 1 7920
box 37576 7920 71256 8880
use CAP_LPF xb36
transform -1 0 37576 0 1 8880
box 37576 8880 71256 9840
use CAP_LPF xb37
transform -1 0 37576 0 1 9840
box 37576 9840 71256 10800
use CAP_LPF xb38
transform -1 0 37576 0 1 10800
box 37576 10800 71256 11760
use CAP_LPF xb39
transform -1 0 37576 0 1 11760
box 37576 11760 71256 12720
use CAP_LPF xb310
transform -1 0 37576 0 1 12720
box 37576 12720 71256 13680
use CAP_LPF xb311
transform -1 0 37576 0 1 13680
box 37576 13680 71256 14640
use CAP_LPF xb312
transform -1 0 37576 0 1 14640
box 37576 14640 71256 15600
use CAP_LPF xb313
transform -1 0 37576 0 1 15600
box 37576 15600 71256 16560
use CAP_LPF xb314
transform -1 0 37576 0 1 16560
box 37576 16560 71256 17520
use CAP_LPF xb315
transform -1 0 37576 0 1 17520
box 37576 17520 71256 18480
use CAP_LPF xb316
transform -1 0 37576 0 1 18480
box 37576 18480 71256 19440
use CAP_LPF xb317
transform -1 0 37576 0 1 19440
box 37576 19440 71256 20400
use CAP_LPF xb318
transform -1 0 37576 0 1 20400
box 37576 20400 71256 21360
use CAP_LPF xb319
transform -1 0 37576 0 1 21360
box 37576 21360 71256 22320
use CAP_LPF xb320
transform -1 0 37576 0 1 22320
box 37576 22320 71256 23280
use CAP_LPF xb321
transform -1 0 37576 0 1 23280
box 37576 23280 71256 24240
use CAP_LPF xb322
transform -1 0 37576 0 1 24240
box 37576 24240 71256 25200
use CAP_LPF xb323
transform -1 0 37576 0 1 25200
box 37576 25200 71256 26160
use cut_M1M4_2x1 
transform 1 0 20596 0 1 0
box 20596 0 20796 76
use cut_M1M2_2x1 
transform 1 0 826 0 1 8122
box 826 8122 1010 8190
use cut_M1M2_2x1 
transform 1 0 2986 0 1 3806
box 2986 3806 3170 3874
use cut_M1M3_2x1 
transform 1 0 826 0 1 12438
box 826 12438 1026 12514
use cut_M1M3_2x1 
transform 1 0 2986 0 1 8122
box 2986 8122 3186 8198
use cut_M1M2_2x1 
transform 1 0 826 0 1 16754
box 826 16754 1010 16822
use cut_M1M2_2x1 
transform 1 0 2986 0 1 12438
box 2986 12438 3170 12506
use cut_M1M3_2x1 
transform 1 0 826 0 1 21070
box 826 21070 1026 21146
use cut_M1M3_2x1 
transform 1 0 2986 0 1 16754
box 2986 16754 3186 16830
use cut_M1M2_2x1 
transform 1 0 2986 0 1 21070
box 2986 21070 3170 21138
use cut_M2M4_2x1 
transform 1 0 3936 0 1 3880
box 3936 3880 4136 3956
use cut_M2M4_2x1 
transform 1 0 3936 0 1 4840
box 3936 4840 4136 4916
use cut_M2M4_2x1 
transform 1 0 3936 0 1 5800
box 3936 5800 4136 5876
use cut_M2M4_2x1 
transform 1 0 3936 0 1 6760
box 3936 6760 4136 6836
use cut_M2M4_2x1 
transform 1 0 3936 0 1 7720
box 3936 7720 4136 7796
use cut_M2M4_2x1 
transform 1 0 3936 0 1 8680
box 3936 8680 4136 8756
use cut_M2M4_2x1 
transform 1 0 3936 0 1 9640
box 3936 9640 4136 9716
use cut_M2M4_2x1 
transform 1 0 3936 0 1 10600
box 3936 10600 4136 10676
use cut_M2M4_2x1 
transform 1 0 3936 0 1 11560
box 3936 11560 4136 11636
use cut_M2M4_2x1 
transform 1 0 3936 0 1 12520
box 3936 12520 4136 12596
use cut_M2M4_2x1 
transform 1 0 3936 0 1 13480
box 3936 13480 4136 13556
use cut_M2M4_2x1 
transform 1 0 3936 0 1 14440
box 3936 14440 4136 14516
use cut_M2M4_2x1 
transform 1 0 3936 0 1 15400
box 3936 15400 4136 15476
use cut_M2M4_2x1 
transform 1 0 3936 0 1 16360
box 3936 16360 4136 16436
use cut_M2M4_2x1 
transform 1 0 3936 0 1 17320
box 3936 17320 4136 17396
use cut_M2M4_2x1 
transform 1 0 3936 0 1 18280
box 3936 18280 4136 18356
use cut_M2M4_2x1 
transform 1 0 3936 0 1 19240
box 3936 19240 4136 19316
use cut_M2M4_2x1 
transform 1 0 3936 0 1 20200
box 3936 20200 4136 20276
use cut_M2M4_2x1 
transform 1 0 3936 0 1 21160
box 3936 21160 4136 21236
use cut_M2M4_2x1 
transform 1 0 3936 0 1 22120
box 3936 22120 4136 22196
use cut_M2M4_2x1 
transform 1 0 3936 0 1 23080
box 3936 23080 4136 23156
use cut_M2M4_2x1 
transform 1 0 3936 0 1 24040
box 3936 24040 4136 24116
use cut_M2M4_2x1 
transform 1 0 3936 0 1 25000
box 3936 25000 4136 25076
use cut_M2M4_2x1 
transform 1 0 3936 0 1 25960
box 3936 25960 4136 26036
use cut_M1M3_2x1 
transform 1 0 826 0 1 3806
box 826 3806 1026 3882
use cut_M3M4_2x1 
transform 1 0 3936 0 1 1000
box 3936 1000 4136 1076
use cut_M3M4_2x1 
transform 1 0 3936 0 1 1960
box 3936 1960 4136 2036
use cut_M3M4_2x1 
transform 1 0 3936 0 1 2920
box 3936 2920 4136 2996
<< labels >>
flabel locali s 37576 0 37816 26400 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 2986 21070 3310 21290 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew
flabel locali s 826 3806 1150 4026 0 FreeSans 400 0 0 0 VLPF
port 3 nsew
<< end >>
