magic
tech sky130A
magscale 1 2
timestamp 1660233442
<< checkpaint >>
rect 112 0 11844 27900
<< m1 >>
rect 2100 10580 2160 27840
rect 2100 10580 2160 27840
rect 1920 140 1980 27840
rect 1920 140 1980 27840
rect 1740 21020 1800 27840
rect 1740 21020 1800 27840
rect 1560 3620 1620 27840
rect 1560 3620 1620 27840
rect 1380 7712 1440 27840
rect 1380 7712 1440 27840
rect 1200 18152 1260 27840
rect 1200 18152 1260 27840
rect 1020 17540 1080 27840
rect 1020 17540 1080 27840
rect 840 19376 900 27840
rect 840 19376 900 27840
rect 660 8936 720 27840
rect 660 8936 720 27840
rect 480 9548 540 27840
rect 480 9548 540 27840
rect 300 8324 360 27840
rect 300 8324 360 27840
rect 120 10160 180 27840
rect 120 10160 180 27840
rect 2668 0 11768 76
<< m2 >>
rect 2160 10642 2340 10718
rect 2160 13702 2340 13778
rect 2160 11866 2340 11942
rect 2160 13090 2340 13166
rect 2160 12478 2340 12554
rect 2160 11254 2340 11330
rect 2160 10642 2340 10718
rect 2160 13702 2340 13778
rect 2160 11866 2340 11942
rect 2160 13090 2340 13166
rect 2160 12478 2340 12554
rect 2160 11254 2340 11330
rect 2160 10642 2340 10718
rect 2160 13702 2340 13778
rect 2160 11866 2340 11942
rect 2160 13090 2340 13166
rect 2160 12478 2340 12554
rect 2160 11254 2340 11330
rect 2160 10642 2340 10718
rect 2160 13702 2340 13778
rect 2160 11866 2340 11942
rect 2160 13090 2340 13166
rect 2160 12478 2340 12554
rect 2160 11254 2340 11330
rect 2160 10642 2340 10718
rect 2160 13702 2340 13778
rect 2160 11866 2340 11942
rect 2160 13090 2340 13166
rect 2160 12478 2340 12554
rect 2160 11254 2340 11330
rect 2160 10642 2340 10718
rect 2160 13702 2340 13778
rect 2160 11866 2340 11942
rect 2160 13090 2340 13166
rect 2160 12478 2340 12554
rect 2160 11254 2340 11330
rect 2160 24562 2340 24638
rect 2160 27622 2340 27698
rect 2160 25786 2340 25862
rect 2160 27010 2340 27086
rect 2160 26398 2340 26474
rect 2160 25174 2340 25250
rect 2160 24562 2340 24638
rect 2160 27622 2340 27698
rect 2160 25786 2340 25862
rect 2160 27010 2340 27086
rect 2160 26398 2340 26474
rect 2160 25174 2340 25250
rect 2160 24562 2340 24638
rect 2160 27622 2340 27698
rect 2160 25786 2340 25862
rect 2160 27010 2340 27086
rect 2160 26398 2340 26474
rect 2160 25174 2340 25250
rect 2160 24562 2340 24638
rect 2160 27622 2340 27698
rect 2160 25786 2340 25862
rect 2160 27010 2340 27086
rect 2160 26398 2340 26474
rect 2160 25174 2340 25250
rect 2160 24562 2340 24638
rect 2160 27622 2340 27698
rect 2160 25786 2340 25862
rect 2160 27010 2340 27086
rect 2160 26398 2340 26474
rect 2160 25174 2340 25250
rect 2160 24562 2340 24638
rect 2160 27622 2340 27698
rect 2160 25786 2340 25862
rect 2160 27010 2340 27086
rect 2160 26398 2340 26474
rect 2160 25174 2340 25250
rect 1980 202 2340 278
rect 1980 3262 2340 3338
rect 1980 1426 2340 1502
rect 1980 2650 2340 2726
rect 1980 2038 2340 2114
rect 1980 814 2340 890
rect 1980 202 2340 278
rect 1980 3262 2340 3338
rect 1980 1426 2340 1502
rect 1980 2650 2340 2726
rect 1980 2038 2340 2114
rect 1980 814 2340 890
rect 1980 202 2340 278
rect 1980 3262 2340 3338
rect 1980 1426 2340 1502
rect 1980 2650 2340 2726
rect 1980 2038 2340 2114
rect 1980 814 2340 890
rect 1980 202 2340 278
rect 1980 3262 2340 3338
rect 1980 1426 2340 1502
rect 1980 2650 2340 2726
rect 1980 2038 2340 2114
rect 1980 814 2340 890
rect 1980 202 2340 278
rect 1980 3262 2340 3338
rect 1980 1426 2340 1502
rect 1980 2650 2340 2726
rect 1980 2038 2340 2114
rect 1980 814 2340 890
rect 1980 202 2340 278
rect 1980 3262 2340 3338
rect 1980 1426 2340 1502
rect 1980 2650 2340 2726
rect 1980 2038 2340 2114
rect 1980 814 2340 890
rect 1980 14122 2340 14198
rect 1980 17182 2340 17258
rect 1980 15346 2340 15422
rect 1980 16570 2340 16646
rect 1980 15958 2340 16034
rect 1980 14734 2340 14810
rect 1980 14122 2340 14198
rect 1980 17182 2340 17258
rect 1980 15346 2340 15422
rect 1980 16570 2340 16646
rect 1980 15958 2340 16034
rect 1980 14734 2340 14810
rect 1980 14122 2340 14198
rect 1980 17182 2340 17258
rect 1980 15346 2340 15422
rect 1980 16570 2340 16646
rect 1980 15958 2340 16034
rect 1980 14734 2340 14810
rect 1980 14122 2340 14198
rect 1980 17182 2340 17258
rect 1980 15346 2340 15422
rect 1980 16570 2340 16646
rect 1980 15958 2340 16034
rect 1980 14734 2340 14810
rect 1980 14122 2340 14198
rect 1980 17182 2340 17258
rect 1980 15346 2340 15422
rect 1980 16570 2340 16646
rect 1980 15958 2340 16034
rect 1980 14734 2340 14810
rect 1980 14122 2340 14198
rect 1980 17182 2340 17258
rect 1980 15346 2340 15422
rect 1980 16570 2340 16646
rect 1980 15958 2340 16034
rect 1980 14734 2340 14810
rect 1800 21082 2340 21158
rect 1800 24142 2340 24218
rect 1800 22306 2340 22382
rect 1800 23530 2340 23606
rect 1800 22918 2340 22994
rect 1800 21694 2340 21770
rect 1800 21082 2340 21158
rect 1800 24142 2340 24218
rect 1800 22306 2340 22382
rect 1800 23530 2340 23606
rect 1800 22918 2340 22994
rect 1800 21694 2340 21770
rect 1800 21082 2340 21158
rect 1800 24142 2340 24218
rect 1800 22306 2340 22382
rect 1800 23530 2340 23606
rect 1800 22918 2340 22994
rect 1800 21694 2340 21770
rect 1800 21082 2340 21158
rect 1800 24142 2340 24218
rect 1800 22306 2340 22382
rect 1800 23530 2340 23606
rect 1800 22918 2340 22994
rect 1800 21694 2340 21770
rect 1800 21082 2340 21158
rect 1800 24142 2340 24218
rect 1800 22306 2340 22382
rect 1800 23530 2340 23606
rect 1800 22918 2340 22994
rect 1800 21694 2340 21770
rect 1800 21082 2340 21158
rect 1800 24142 2340 24218
rect 1800 22306 2340 22382
rect 1800 23530 2340 23606
rect 1800 22918 2340 22994
rect 1800 21694 2340 21770
rect 1620 3682 2340 3758
rect 1620 6742 2340 6818
rect 1620 4906 2340 4982
rect 1620 6130 2340 6206
rect 1620 5518 2340 5594
rect 1620 4294 2340 4370
rect 1620 3682 2340 3758
rect 1620 6742 2340 6818
rect 1620 4906 2340 4982
rect 1620 6130 2340 6206
rect 1620 5518 2340 5594
rect 1620 4294 2340 4370
rect 1620 3682 2340 3758
rect 1620 6742 2340 6818
rect 1620 4906 2340 4982
rect 1620 6130 2340 6206
rect 1620 5518 2340 5594
rect 1620 4294 2340 4370
rect 1620 3682 2340 3758
rect 1620 6742 2340 6818
rect 1620 4906 2340 4982
rect 1620 6130 2340 6206
rect 1620 5518 2340 5594
rect 1620 4294 2340 4370
rect 1620 3682 2340 3758
rect 1620 6742 2340 6818
rect 1620 4906 2340 4982
rect 1620 6130 2340 6206
rect 1620 5518 2340 5594
rect 1620 4294 2340 4370
rect 1620 3682 2340 3758
rect 1620 6742 2340 6818
rect 1620 4906 2340 4982
rect 1620 6130 2340 6206
rect 1620 5518 2340 5594
rect 1620 4294 2340 4370
rect 1440 7774 2340 7850
rect 1260 18214 2340 18290
rect 1080 17602 2340 17678
rect 1080 20662 2340 20738
rect 1080 18826 2340 18902
rect 1080 20050 2340 20126
rect 1080 17602 2340 17678
rect 1080 20662 2340 20738
rect 1080 18826 2340 18902
rect 1080 20050 2340 20126
rect 1080 17602 2340 17678
rect 1080 20662 2340 20738
rect 1080 18826 2340 18902
rect 1080 20050 2340 20126
rect 1080 17602 2340 17678
rect 1080 20662 2340 20738
rect 1080 18826 2340 18902
rect 1080 20050 2340 20126
rect 900 19438 2340 19514
rect 720 8998 2340 9074
rect 540 9610 2340 9686
rect 360 8386 2340 8462
rect 180 10222 2340 10298
<< m3 >>
rect 2668 24360 2744 27900
use SUNSAR_CAP32C_CV XC1
transform 1 0 2340 0 1 0
box 2340 0 11844 3480
use SUNSAR_CAP32C_CV XC64a<0>
transform 1 0 2340 0 1 3480
box 2340 3480 11844 6960
use SUNSAR_CAP32C_CV XC32a<0>
transform 1 0 2340 0 1 6960
box 2340 6960 11844 10440
use SUNSAR_CAP32C_CV XC128a<1>
transform 1 0 2340 0 1 10440
box 2340 10440 11844 13920
use SUNSAR_CAP32C_CV XC128b<2>
transform 1 0 2340 0 1 13920
box 2340 13920 11844 17400
use SUNSAR_CAP32C_CV X16ab
transform 1 0 2340 0 1 17400
box 2340 17400 11844 20880
use SUNSAR_CAP32C_CV XC64b<1>
transform 1 0 2340 0 1 20880
box 2340 20880 11844 24360
use SUNSAR_CAP32C_CV XC0
transform 1 0 2340 0 1 24360
box 2340 24360 11844 27840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10642
box 2340 10642 2540 10718
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 10580
box 2092 10580 2168 10780
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13702
box 2340 13702 2540 13778
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13640
box 2092 13640 2168 13840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11866
box 2340 11866 2540 11942
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11804
box 2092 11804 2168 12004
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13090
box 2340 13090 2540 13166
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13028
box 2092 13028 2168 13228
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 12478
box 2340 12478 2540 12554
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 12416
box 2092 12416 2168 12616
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11254
box 2340 11254 2540 11330
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11192
box 2092 11192 2168 11392
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10642
box 2340 10642 2540 10718
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 10580
box 2092 10580 2168 10780
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13702
box 2340 13702 2540 13778
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13640
box 2092 13640 2168 13840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11866
box 2340 11866 2540 11942
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11804
box 2092 11804 2168 12004
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13090
box 2340 13090 2540 13166
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13028
box 2092 13028 2168 13228
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 12478
box 2340 12478 2540 12554
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 12416
box 2092 12416 2168 12616
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11254
box 2340 11254 2540 11330
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11192
box 2092 11192 2168 11392
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10642
box 2340 10642 2540 10718
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 10580
box 2092 10580 2168 10780
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13702
box 2340 13702 2540 13778
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13640
box 2092 13640 2168 13840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11866
box 2340 11866 2540 11942
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11804
box 2092 11804 2168 12004
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13090
box 2340 13090 2540 13166
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13028
box 2092 13028 2168 13228
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 12478
box 2340 12478 2540 12554
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 12416
box 2092 12416 2168 12616
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11254
box 2340 11254 2540 11330
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11192
box 2092 11192 2168 11392
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10642
box 2340 10642 2540 10718
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 10580
box 2092 10580 2168 10780
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13702
box 2340 13702 2540 13778
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13640
box 2092 13640 2168 13840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11866
box 2340 11866 2540 11942
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11804
box 2092 11804 2168 12004
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13090
box 2340 13090 2540 13166
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13028
box 2092 13028 2168 13228
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 12478
box 2340 12478 2540 12554
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 12416
box 2092 12416 2168 12616
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11254
box 2340 11254 2540 11330
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11192
box 2092 11192 2168 11392
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10642
box 2340 10642 2540 10718
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 10580
box 2092 10580 2168 10780
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13702
box 2340 13702 2540 13778
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13640
box 2092 13640 2168 13840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11866
box 2340 11866 2540 11942
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11804
box 2092 11804 2168 12004
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13090
box 2340 13090 2540 13166
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13028
box 2092 13028 2168 13228
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 12478
box 2340 12478 2540 12554
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 12416
box 2092 12416 2168 12616
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11254
box 2340 11254 2540 11330
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11192
box 2092 11192 2168 11392
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10642
box 2340 10642 2540 10718
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 10580
box 2092 10580 2168 10780
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13702
box 2340 13702 2540 13778
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13640
box 2092 13640 2168 13840
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11866
box 2340 11866 2540 11942
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11804
box 2092 11804 2168 12004
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 13090
box 2340 13090 2540 13166
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 13028
box 2092 13028 2168 13228
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 12478
box 2340 12478 2540 12554
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 12416
box 2092 12416 2168 12616
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 11254
box 2340 11254 2540 11330
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 11192
box 2092 11192 2168 11392
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24562
box 2340 24562 2540 24638
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 24500
box 2092 24500 2168 24700
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27622
box 2340 27622 2540 27698
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 27560
box 2092 27560 2168 27760
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25786
box 2340 25786 2540 25862
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25724
box 2092 25724 2168 25924
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27010
box 2340 27010 2540 27086
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26948
box 2092 26948 2168 27148
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 26398
box 2340 26398 2540 26474
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26336
box 2092 26336 2168 26536
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25174
box 2340 25174 2540 25250
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25112
box 2092 25112 2168 25312
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24562
box 2340 24562 2540 24638
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 24500
box 2092 24500 2168 24700
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27622
box 2340 27622 2540 27698
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 27560
box 2092 27560 2168 27760
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25786
box 2340 25786 2540 25862
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25724
box 2092 25724 2168 25924
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27010
box 2340 27010 2540 27086
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26948
box 2092 26948 2168 27148
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 26398
box 2340 26398 2540 26474
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26336
box 2092 26336 2168 26536
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25174
box 2340 25174 2540 25250
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25112
box 2092 25112 2168 25312
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24562
box 2340 24562 2540 24638
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 24500
box 2092 24500 2168 24700
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27622
box 2340 27622 2540 27698
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 27560
box 2092 27560 2168 27760
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25786
box 2340 25786 2540 25862
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25724
box 2092 25724 2168 25924
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27010
box 2340 27010 2540 27086
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26948
box 2092 26948 2168 27148
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 26398
box 2340 26398 2540 26474
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26336
box 2092 26336 2168 26536
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25174
box 2340 25174 2540 25250
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25112
box 2092 25112 2168 25312
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24562
box 2340 24562 2540 24638
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 24500
box 2092 24500 2168 24700
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27622
box 2340 27622 2540 27698
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 27560
box 2092 27560 2168 27760
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25786
box 2340 25786 2540 25862
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25724
box 2092 25724 2168 25924
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27010
box 2340 27010 2540 27086
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26948
box 2092 26948 2168 27148
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 26398
box 2340 26398 2540 26474
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26336
box 2092 26336 2168 26536
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25174
box 2340 25174 2540 25250
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25112
box 2092 25112 2168 25312
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24562
box 2340 24562 2540 24638
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 24500
box 2092 24500 2168 24700
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27622
box 2340 27622 2540 27698
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 27560
box 2092 27560 2168 27760
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25786
box 2340 25786 2540 25862
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25724
box 2092 25724 2168 25924
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27010
box 2340 27010 2540 27086
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26948
box 2092 26948 2168 27148
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 26398
box 2340 26398 2540 26474
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26336
box 2092 26336 2168 26536
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25174
box 2340 25174 2540 25250
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25112
box 2092 25112 2168 25312
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24562
box 2340 24562 2540 24638
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 24500
box 2092 24500 2168 24700
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27622
box 2340 27622 2540 27698
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 27560
box 2092 27560 2168 27760
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25786
box 2340 25786 2540 25862
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25724
box 2092 25724 2168 25924
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 27010
box 2340 27010 2540 27086
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26948
box 2092 26948 2168 27148
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 26398
box 2340 26398 2540 26474
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 26336
box 2092 26336 2168 26536
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 25174
box 2340 25174 2540 25250
use SUNSAR_cut_M2M3_1x2 
transform 1 0 2092 0 1 25112
box 2092 25112 2168 25312
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3262
box 2340 3262 2540 3338
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 3200
box 1912 3200 1988 3400
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 1426
box 2340 1426 2540 1502
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1364
box 1912 1364 1988 1564
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2650
box 2340 2650 2540 2726
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 2588
box 1912 2588 1988 2788
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2038
box 2340 2038 2540 2114
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1976
box 1912 1976 1988 2176
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 814
box 2340 814 2540 890
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 752
box 1912 752 1988 952
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3262
box 2340 3262 2540 3338
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 3200
box 1912 3200 1988 3400
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 1426
box 2340 1426 2540 1502
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1364
box 1912 1364 1988 1564
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2650
box 2340 2650 2540 2726
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 2588
box 1912 2588 1988 2788
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2038
box 2340 2038 2540 2114
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1976
box 1912 1976 1988 2176
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 814
box 2340 814 2540 890
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 752
box 1912 752 1988 952
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3262
box 2340 3262 2540 3338
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 3200
box 1912 3200 1988 3400
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 1426
box 2340 1426 2540 1502
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1364
box 1912 1364 1988 1564
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2650
box 2340 2650 2540 2726
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 2588
box 1912 2588 1988 2788
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2038
box 2340 2038 2540 2114
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1976
box 1912 1976 1988 2176
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 814
box 2340 814 2540 890
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 752
box 1912 752 1988 952
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3262
box 2340 3262 2540 3338
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 3200
box 1912 3200 1988 3400
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 1426
box 2340 1426 2540 1502
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1364
box 1912 1364 1988 1564
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2650
box 2340 2650 2540 2726
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 2588
box 1912 2588 1988 2788
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2038
box 2340 2038 2540 2114
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1976
box 1912 1976 1988 2176
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 814
box 2340 814 2540 890
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 752
box 1912 752 1988 952
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3262
box 2340 3262 2540 3338
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 3200
box 1912 3200 1988 3400
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 1426
box 2340 1426 2540 1502
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1364
box 1912 1364 1988 1564
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2650
box 2340 2650 2540 2726
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 2588
box 1912 2588 1988 2788
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2038
box 2340 2038 2540 2114
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1976
box 1912 1976 1988 2176
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 814
box 2340 814 2540 890
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 752
box 1912 752 1988 952
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3262
box 2340 3262 2540 3338
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 3200
box 1912 3200 1988 3400
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 1426
box 2340 1426 2540 1502
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1364
box 1912 1364 1988 1564
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2650
box 2340 2650 2540 2726
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 2588
box 1912 2588 1988 2788
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 2038
box 2340 2038 2540 2114
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 1976
box 1912 1976 1988 2176
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 814
box 2340 814 2540 890
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 752
box 1912 752 1988 952
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14122
box 2340 14122 2540 14198
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14060
box 1912 14060 1988 14260
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17182
box 2340 17182 2540 17258
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 17120
box 1912 17120 1988 17320
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15346
box 2340 15346 2540 15422
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15284
box 1912 15284 1988 15484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 16570
box 2340 16570 2540 16646
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 16508
box 1912 16508 1988 16708
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15958
box 2340 15958 2540 16034
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15896
box 1912 15896 1988 16096
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14734
box 2340 14734 2540 14810
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14672
box 1912 14672 1988 14872
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14122
box 2340 14122 2540 14198
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14060
box 1912 14060 1988 14260
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17182
box 2340 17182 2540 17258
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 17120
box 1912 17120 1988 17320
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15346
box 2340 15346 2540 15422
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15284
box 1912 15284 1988 15484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 16570
box 2340 16570 2540 16646
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 16508
box 1912 16508 1988 16708
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15958
box 2340 15958 2540 16034
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15896
box 1912 15896 1988 16096
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14734
box 2340 14734 2540 14810
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14672
box 1912 14672 1988 14872
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14122
box 2340 14122 2540 14198
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14060
box 1912 14060 1988 14260
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17182
box 2340 17182 2540 17258
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 17120
box 1912 17120 1988 17320
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15346
box 2340 15346 2540 15422
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15284
box 1912 15284 1988 15484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 16570
box 2340 16570 2540 16646
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 16508
box 1912 16508 1988 16708
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15958
box 2340 15958 2540 16034
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15896
box 1912 15896 1988 16096
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14734
box 2340 14734 2540 14810
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14672
box 1912 14672 1988 14872
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14122
box 2340 14122 2540 14198
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14060
box 1912 14060 1988 14260
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17182
box 2340 17182 2540 17258
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 17120
box 1912 17120 1988 17320
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15346
box 2340 15346 2540 15422
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15284
box 1912 15284 1988 15484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 16570
box 2340 16570 2540 16646
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 16508
box 1912 16508 1988 16708
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15958
box 2340 15958 2540 16034
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15896
box 1912 15896 1988 16096
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14734
box 2340 14734 2540 14810
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14672
box 1912 14672 1988 14872
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14122
box 2340 14122 2540 14198
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14060
box 1912 14060 1988 14260
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17182
box 2340 17182 2540 17258
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 17120
box 1912 17120 1988 17320
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15346
box 2340 15346 2540 15422
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15284
box 1912 15284 1988 15484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 16570
box 2340 16570 2540 16646
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 16508
box 1912 16508 1988 16708
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15958
box 2340 15958 2540 16034
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15896
box 1912 15896 1988 16096
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14734
box 2340 14734 2540 14810
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14672
box 1912 14672 1988 14872
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14122
box 2340 14122 2540 14198
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14060
box 1912 14060 1988 14260
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17182
box 2340 17182 2540 17258
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 17120
box 1912 17120 1988 17320
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15346
box 2340 15346 2540 15422
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15284
box 1912 15284 1988 15484
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 16570
box 2340 16570 2540 16646
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 16508
box 1912 16508 1988 16708
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 15958
box 2340 15958 2540 16034
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 15896
box 1912 15896 1988 16096
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 14734
box 2340 14734 2540 14810
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1912 0 1 14672
box 1912 14672 1988 14872
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21082
box 2340 21082 2540 21158
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21020
box 1732 21020 1808 21220
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24142
box 2340 24142 2540 24218
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 24080
box 1732 24080 1808 24280
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22306
box 2340 22306 2540 22382
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22244
box 1732 22244 1808 22444
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 23530
box 2340 23530 2540 23606
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 23468
box 1732 23468 1808 23668
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22918
box 2340 22918 2540 22994
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22856
box 1732 22856 1808 23056
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21694
box 2340 21694 2540 21770
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21632
box 1732 21632 1808 21832
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21082
box 2340 21082 2540 21158
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21020
box 1732 21020 1808 21220
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24142
box 2340 24142 2540 24218
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 24080
box 1732 24080 1808 24280
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22306
box 2340 22306 2540 22382
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22244
box 1732 22244 1808 22444
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 23530
box 2340 23530 2540 23606
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 23468
box 1732 23468 1808 23668
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22918
box 2340 22918 2540 22994
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22856
box 1732 22856 1808 23056
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21694
box 2340 21694 2540 21770
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21632
box 1732 21632 1808 21832
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21082
box 2340 21082 2540 21158
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21020
box 1732 21020 1808 21220
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24142
box 2340 24142 2540 24218
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 24080
box 1732 24080 1808 24280
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22306
box 2340 22306 2540 22382
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22244
box 1732 22244 1808 22444
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 23530
box 2340 23530 2540 23606
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 23468
box 1732 23468 1808 23668
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22918
box 2340 22918 2540 22994
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22856
box 1732 22856 1808 23056
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21694
box 2340 21694 2540 21770
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21632
box 1732 21632 1808 21832
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21082
box 2340 21082 2540 21158
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21020
box 1732 21020 1808 21220
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24142
box 2340 24142 2540 24218
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 24080
box 1732 24080 1808 24280
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22306
box 2340 22306 2540 22382
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22244
box 1732 22244 1808 22444
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 23530
box 2340 23530 2540 23606
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 23468
box 1732 23468 1808 23668
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22918
box 2340 22918 2540 22994
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22856
box 1732 22856 1808 23056
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21694
box 2340 21694 2540 21770
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21632
box 1732 21632 1808 21832
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21082
box 2340 21082 2540 21158
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21020
box 1732 21020 1808 21220
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24142
box 2340 24142 2540 24218
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 24080
box 1732 24080 1808 24280
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22306
box 2340 22306 2540 22382
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22244
box 1732 22244 1808 22444
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 23530
box 2340 23530 2540 23606
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 23468
box 1732 23468 1808 23668
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22918
box 2340 22918 2540 22994
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22856
box 1732 22856 1808 23056
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21694
box 2340 21694 2540 21770
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21632
box 1732 21632 1808 21832
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21082
box 2340 21082 2540 21158
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21020
box 1732 21020 1808 21220
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 24142
box 2340 24142 2540 24218
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 24080
box 1732 24080 1808 24280
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22306
box 2340 22306 2540 22382
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22244
box 1732 22244 1808 22444
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 23530
box 2340 23530 2540 23606
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 23468
box 1732 23468 1808 23668
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 22918
box 2340 22918 2540 22994
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 22856
box 1732 22856 1808 23056
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 21694
box 2340 21694 2540 21770
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1732 0 1 21632
box 1732 21632 1808 21832
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3682
box 2340 3682 2540 3758
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 3620
box 1552 3620 1628 3820
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6742
box 2340 6742 2540 6818
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6680
box 1552 6680 1628 6880
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4906
box 2340 4906 2540 4982
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4844
box 1552 4844 1628 5044
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6130
box 2340 6130 2540 6206
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6068
box 1552 6068 1628 6268
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 5518
box 2340 5518 2540 5594
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 5456
box 1552 5456 1628 5656
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4294
box 2340 4294 2540 4370
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4232
box 1552 4232 1628 4432
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3682
box 2340 3682 2540 3758
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 3620
box 1552 3620 1628 3820
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6742
box 2340 6742 2540 6818
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6680
box 1552 6680 1628 6880
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4906
box 2340 4906 2540 4982
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4844
box 1552 4844 1628 5044
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6130
box 2340 6130 2540 6206
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6068
box 1552 6068 1628 6268
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 5518
box 2340 5518 2540 5594
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 5456
box 1552 5456 1628 5656
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4294
box 2340 4294 2540 4370
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4232
box 1552 4232 1628 4432
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3682
box 2340 3682 2540 3758
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 3620
box 1552 3620 1628 3820
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6742
box 2340 6742 2540 6818
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6680
box 1552 6680 1628 6880
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4906
box 2340 4906 2540 4982
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4844
box 1552 4844 1628 5044
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6130
box 2340 6130 2540 6206
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6068
box 1552 6068 1628 6268
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 5518
box 2340 5518 2540 5594
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 5456
box 1552 5456 1628 5656
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4294
box 2340 4294 2540 4370
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4232
box 1552 4232 1628 4432
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3682
box 2340 3682 2540 3758
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 3620
box 1552 3620 1628 3820
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6742
box 2340 6742 2540 6818
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6680
box 1552 6680 1628 6880
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4906
box 2340 4906 2540 4982
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4844
box 1552 4844 1628 5044
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6130
box 2340 6130 2540 6206
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6068
box 1552 6068 1628 6268
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 5518
box 2340 5518 2540 5594
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 5456
box 1552 5456 1628 5656
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4294
box 2340 4294 2540 4370
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4232
box 1552 4232 1628 4432
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3682
box 2340 3682 2540 3758
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 3620
box 1552 3620 1628 3820
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6742
box 2340 6742 2540 6818
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6680
box 1552 6680 1628 6880
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4906
box 2340 4906 2540 4982
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4844
box 1552 4844 1628 5044
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6130
box 2340 6130 2540 6206
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6068
box 1552 6068 1628 6268
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 5518
box 2340 5518 2540 5594
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 5456
box 1552 5456 1628 5656
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4294
box 2340 4294 2540 4370
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4232
box 1552 4232 1628 4432
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 3682
box 2340 3682 2540 3758
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 3620
box 1552 3620 1628 3820
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6742
box 2340 6742 2540 6818
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6680
box 1552 6680 1628 6880
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4906
box 2340 4906 2540 4982
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4844
box 1552 4844 1628 5044
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 6130
box 2340 6130 2540 6206
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 6068
box 1552 6068 1628 6268
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 5518
box 2340 5518 2540 5594
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 5456
box 1552 5456 1628 5656
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 4294
box 2340 4294 2540 4370
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1552 0 1 4232
box 1552 4232 1628 4432
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 7774
box 2340 7774 2540 7850
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1372 0 1 7712
box 1372 7712 1448 7912
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 18214
box 2340 18214 2540 18290
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1192 0 1 18152
box 1192 18152 1268 18352
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17602
box 2340 17602 2540 17678
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 17540
box 1012 17540 1088 17740
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20662
box 2340 20662 2540 20738
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 20600
box 1012 20600 1088 20800
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 18826
box 2340 18826 2540 18902
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 18764
box 1012 18764 1088 18964
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20050
box 2340 20050 2540 20126
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 19988
box 1012 19988 1088 20188
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17602
box 2340 17602 2540 17678
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 17540
box 1012 17540 1088 17740
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20662
box 2340 20662 2540 20738
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 20600
box 1012 20600 1088 20800
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 18826
box 2340 18826 2540 18902
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 18764
box 1012 18764 1088 18964
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20050
box 2340 20050 2540 20126
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 19988
box 1012 19988 1088 20188
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17602
box 2340 17602 2540 17678
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 17540
box 1012 17540 1088 17740
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20662
box 2340 20662 2540 20738
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 20600
box 1012 20600 1088 20800
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 18826
box 2340 18826 2540 18902
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 18764
box 1012 18764 1088 18964
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20050
box 2340 20050 2540 20126
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 19988
box 1012 19988 1088 20188
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 17602
box 2340 17602 2540 17678
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 17540
box 1012 17540 1088 17740
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20662
box 2340 20662 2540 20738
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 20600
box 1012 20600 1088 20800
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 18826
box 2340 18826 2540 18902
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 18764
box 1012 18764 1088 18964
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 20050
box 2340 20050 2540 20126
use SUNSAR_cut_M2M3_1x2 
transform 1 0 1012 0 1 19988
box 1012 19988 1088 20188
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 19438
box 2340 19438 2540 19514
use SUNSAR_cut_M2M3_1x2 
transform 1 0 832 0 1 19376
box 832 19376 908 19576
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 8998
box 2340 8998 2540 9074
use SUNSAR_cut_M2M3_1x2 
transform 1 0 652 0 1 8936
box 652 8936 728 9136
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 9610
box 2340 9610 2540 9686
use SUNSAR_cut_M2M3_1x2 
transform 1 0 472 0 1 9548
box 472 9548 548 9748
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 8386
box 2340 8386 2540 8462
use SUNSAR_cut_M2M3_1x2 
transform 1 0 292 0 1 8324
box 292 8324 368 8524
use SUNSAR_cut_M1M3_2x1 
transform 1 0 2340 0 1 10222
box 2340 10222 2540 10298
use SUNSAR_cut_M2M3_1x2 
transform 1 0 112 0 1 10160
box 112 10160 188 10360
use SUNSAR_cut_M1M2_1x2 
transform 1 0 2668 0 1 7108
box 2668 7108 2736 7292
use SUNSAR_cut_M1M2_1x2 
transform 1 0 2668 0 1 7108
box 2668 7108 2736 7292
<< labels >>
flabel m1 s 2100 10580 2160 27840 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew
flabel m1 s 1920 140 1980 27840 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew
flabel m1 s 1740 21020 1800 27840 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew
flabel m1 s 1560 3620 1620 27840 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew
flabel m1 s 1380 7712 1440 27840 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew
flabel m1 s 1200 18152 1260 27840 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew
flabel m1 s 1020 17540 1080 27840 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew
flabel m1 s 840 19376 900 27840 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew
flabel m1 s 660 8936 720 27840 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew
flabel m1 s 480 9548 540 27840 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew
flabel m1 s 300 8324 360 27840 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew
flabel m1 s 120 10160 180 27840 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew
flabel m1 s 2668 0 11768 76 0 FreeSans 400 0 0 0 AVSS
port 14 nsew
flabel m3 s 2668 24360 2744 27900 0 FreeSans 400 0 0 0 CTOP
port 13 nsew
<< end >>
