magic
tech sky130A
magscale 1 2
timestamp 1661983200
<< checkpaint >>
rect 0 0 4416 10688
<< locali >>
rect 3792 384 4032 10304
rect 384 384 4032 624
rect 384 10064 4032 10304
rect 384 384 624 10304
rect 3792 384 4032 10304
rect 4176 0 4416 10688
rect 0 0 4416 240
rect 0 10448 4416 10688
rect 0 0 240 10688
rect 4176 0 4416 10688
rect 1200 4786 1368 4846
rect 1200 5314 1368 5374
rect 1200 5842 1368 5902
rect 1200 6370 1368 6430
rect 1200 6898 1368 6958
rect 1200 7426 1368 7486
rect 1200 7954 1368 8014
rect 1200 8482 1368 8542
rect 1200 9010 1368 9070
rect 1200 9538 1368 9598
rect 1368 4786 1428 9598
rect 3252 1706 3420 1766
rect 3252 1882 3420 1942
rect 3420 1706 3480 1942
rect 1170 914 1230 2734
rect 1632 4170 1800 4230
rect 1632 4346 1800 4406
rect 1800 4170 1860 4406
rect 1632 826 2004 886
rect 1632 2586 2004 2646
rect 2004 826 2064 2646
rect 1632 826 2004 886
rect 1632 4698 2004 4758
rect 1632 5226 2004 5286
rect 1632 5754 2004 5814
rect 1632 6282 2004 6342
rect 1632 6810 2004 6870
rect 1632 7338 2004 7398
rect 1632 7866 2004 7926
rect 1632 8394 2004 8454
rect 1632 8922 2004 8982
rect 1632 9450 2004 9510
rect 2004 826 2064 9510
rect 3252 826 3624 886
rect 3252 1354 3624 1414
rect 3624 826 3684 1414
rect 3252 826 3624 886
rect 3252 2234 3624 2294
rect 3624 826 3684 2294
<< m1 >>
rect 1524 384 1740 886
rect 660 384 876 988
rect 3144 0 3360 886
rect 2280 0 2496 988
rect 2820 914 2988 974
rect 2988 1178 3252 1238
rect 1632 2410 2988 2470
rect 2820 1442 2988 1502
rect 2988 914 3048 2478
rect 3252 2058 3420 2118
rect 1632 4522 3420 4582
rect 3252 2410 3420 2470
rect 3420 2058 3480 4590
rect 1632 4874 1800 4934
rect 1632 5402 1800 5462
rect 1632 5930 1800 5990
rect 1632 6458 1800 6518
rect 1632 6986 1800 7046
rect 1632 7514 1800 7574
rect 1632 8042 1800 8102
rect 1632 8570 1800 8630
rect 1632 9098 1800 9158
rect 1632 9626 1800 9686
rect 1800 4874 1860 9694
<< m2 >>
rect 0 1970 216 2030
rect 4200 4522 4416 4582
rect 0 4434 216 4494
rect 0 914 216 974
rect 4200 4874 4416 4934
rect 0 2322 216 2382
rect 0 4786 216 4846
rect 0 2322 216 2382
rect 2572 2292 2820 2368
rect 108 2322 2572 2398
rect 2572 2284 2648 2398
rect 0 4786 216 4846
rect 952 4786 1200 4862
rect 108 4786 952 4862
rect 952 4786 1028 4862
rect 0 914 216 974
rect 952 914 1200 990
rect 108 914 952 990
rect 952 914 1028 990
rect 4200 4522 4416 4582
rect 1632 4522 1804 4598
rect 1804 4522 4308 4598
rect 1804 4522 1880 4598
rect 4200 4874 4416 4934
rect 1632 4874 1804 4950
rect 1804 4874 4308 4950
rect 1804 4874 1880 4950
rect 0 1970 216 2030
rect 2572 1970 2820 2046
rect 108 1970 2572 2046
rect 2572 1970 2648 2046
rect 0 4434 216 4494
rect 952 4434 1200 4510
rect 108 4434 952 4510
rect 952 4434 1028 4510
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa10
transform 1 0 768 0 1 768
box 768 768 2028 2528
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa20
transform 1 0 768 0 1 2528
box 768 2528 2028 4288
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa30
transform 1 0 768 0 1 4288
box 768 4288 2028 4640
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa40
transform 1 0 768 0 1 4640
box 768 4640 2028 5168
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa41
transform 1 0 768 0 1 5168
box 768 5168 2028 5696
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa42
transform 1 0 768 0 1 5696
box 768 5696 2028 6224
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa43
transform 1 0 768 0 1 6224
box 768 6224 2028 6752
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa44
transform 1 0 768 0 1 6752
box 768 6752 2028 7280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa45
transform 1 0 768 0 1 7280
box 768 7280 2028 7808
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa46
transform 1 0 768 0 1 7808
box 768 7808 2028 8336
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa47
transform 1 0 768 0 1 8336
box 768 8336 2028 8864
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa48
transform 1 0 768 0 1 8864
box 768 8864 2028 9392
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa49
transform 1 0 768 0 1 9392
box 768 9392 2028 9920
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM xb10
transform -1 0 3648 0 1 768
box 3648 768 4908 1296
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM xb20
transform -1 0 3648 0 1 1296
box 3648 1296 4908 1824
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xb30
transform -1 0 3648 0 1 1824
box 3648 1824 4908 2176
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xb40
transform -1 0 3648 0 1 2176
box 3648 2176 4908 2528
use cut_M1M2_2x1 
transform 1 0 1540 0 1 826
box 1540 826 1724 894
use cut_M1M2_2x1 
transform 1 0 1540 0 1 384
box 1540 384 1724 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 900
box 676 900 860 968
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 3160 0 1 826
box 3160 826 3344 894
use cut_M1M2_2x1 
transform 1 0 3160 0 1 0
box 3160 0 3344 68
use cut_M1M2_2x1 
transform 1 0 2296 0 1 900
box 2296 900 2480 968
use cut_M1M2_2x1 
transform 1 0 2296 0 1 0
box 2296 0 2480 68
use cut_M1M2_2x1 
transform 1 0 2712 0 1 914
box 2712 914 2896 982
use cut_M1M2_2x1 
transform 1 0 3144 0 1 1178
box 3144 1178 3328 1246
use cut_M1M2_2x1 
transform 1 0 1524 0 1 2410
box 1524 2410 1708 2478
use cut_M1M2_2x1 
transform 1 0 2712 0 1 1442
box 2712 1442 2896 1510
use cut_M1M2_2x1 
transform 1 0 3144 0 1 2058
box 3144 2058 3328 2126
use cut_M1M2_2x1 
transform 1 0 1524 0 1 4522
box 1524 4522 1708 4590
use cut_M1M2_2x1 
transform 1 0 3144 0 1 2410
box 3144 2410 3328 2478
use cut_M1M2_2x1 
transform 1 0 1524 0 1 4874
box 1524 4874 1708 4942
use cut_M1M2_2x1 
transform 1 0 1524 0 1 5402
box 1524 5402 1708 5470
use cut_M1M2_2x1 
transform 1 0 1524 0 1 5930
box 1524 5930 1708 5998
use cut_M1M2_2x1 
transform 1 0 1524 0 1 6458
box 1524 6458 1708 6526
use cut_M1M2_2x1 
transform 1 0 1524 0 1 6986
box 1524 6986 1708 7054
use cut_M1M2_2x1 
transform 1 0 1524 0 1 7514
box 1524 7514 1708 7582
use cut_M1M2_2x1 
transform 1 0 1524 0 1 8042
box 1524 8042 1708 8110
use cut_M1M2_2x1 
transform 1 0 1524 0 1 8570
box 1524 8570 1708 8638
use cut_M1M2_2x1 
transform 1 0 1524 0 1 9098
box 1524 9098 1708 9166
use cut_M1M2_2x1 
transform 1 0 1524 0 1 9626
box 1524 9626 1708 9694
use cut_M1M3_2x1 
transform 1 0 2728 0 1 2284
box 2728 2284 2928 2360
use cut_M1M3_2x1 
transform 1 0 1108 0 1 4786
box 1108 4786 1308 4862
use cut_M1M3_2x1 
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M3_2x1 
transform 1 0 1524 0 1 4522
box 1524 4522 1724 4598
use cut_M1M3_2x1 
transform 1 0 1524 0 1 4874
box 1524 4874 1724 4950
use cut_M1M3_2x1 
transform 1 0 2728 0 1 1970
box 2728 1970 2928 2046
use cut_M1M3_2x1 
transform 1 0 1108 0 1 4434
box 1108 4434 1308 4510
<< labels >>
flabel locali s 3792 384 4032 10304 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 4176 0 4416 10688 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 0 1970 216 2030 0 FreeSans 400 0 0 0 CP_UP_N
port 2 nsew
flabel m2 s 4200 4522 4416 4582 0 FreeSans 400 0 0 0 LPF
port 3 nsew
flabel m2 s 0 4434 216 4494 0 FreeSans 400 0 0 0 CP_DOWN
port 4 nsew
flabel m2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew
flabel m2 s 4200 4874 4416 4934 0 FreeSans 400 0 0 0 LPFZ
port 7 nsew
flabel m2 s 0 2322 216 2382 0 FreeSans 400 0 0 0 PWRUP_1V8
port 8 nsew
flabel m2 s 0 4786 216 4846 0 FreeSans 400 0 0 0 KICK
port 9 nsew
<< end >>
