magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 2240
<< poly >>
rect 270 2062 1710 2098
rect 270 142 1710 178
<< locali >>
rect 1590 1410 1650 2110
rect 330 450 390 1790
rect 720 530 858 590
rect 720 1170 858 1230
rect 720 1810 858 1870
rect 858 530 1260 590
rect 858 530 918 1870
rect 522 210 720 270
rect 522 850 720 910
rect 522 1490 720 1550
rect 522 210 582 1550
rect 720 210 858 270
rect 858 50 1260 110
rect 858 50 918 270
rect 1062 1170 1260 1230
rect 1062 1810 1260 1870
rect 720 2130 1062 2190
rect 1062 1170 1122 2190
rect 1620 130 1758 190
rect 1620 450 1758 510
rect 1620 1090 1758 1150
rect 1758 130 1818 1150
rect 690 210 750 430
rect 690 530 750 750
rect 690 850 750 1070
rect 690 1170 750 1390
rect 690 1490 750 1710
rect 690 1810 750 2030
rect 1230 210 1290 430
rect 1230 530 1290 750
rect 1230 850 1290 1070
rect 1230 1170 1290 1390
rect 1230 1490 1290 1710
rect 1230 1810 1290 2030
<< m3 >>
rect 1260 850 1398 910
rect 1398 770 1620 830
rect 1398 770 1458 918
rect 1170 0 1354 2240
rect 630 0 814 2240
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 990 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 990 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 990 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 990 1280
use NCHDL MN4
transform 1 0 0 0 1 1280
box 0 1280 990 1600
use NCHDL MN5
transform 1 0 0 0 1 1600
box 0 1600 990 1920
use NCHDL MN6
transform 1 0 0 0 1 1920
box 0 1920 990 2240
use PCHDL MP0
transform 1 0 990 0 1 0
box 990 0 1980 320
use PCHDL MP1
transform 1 0 990 0 1 320
box 990 320 1980 640
use PCHDL MP2
transform 1 0 990 0 1 640
box 990 640 1980 960
use PCHDL MP3
transform 1 0 990 0 1 960
box 990 960 1980 1280
use PCHDL MP4
transform 1 0 990 0 1 1280
box 990 1280 1980 1600
use PCHDL MP5
transform 1 0 990 0 1 1600
box 990 1600 1980 1920
use PCHDL MP6
transform 1 0 990 0 1 1920
box 990 1920 1980 2240
use cut_M1M4_2x1 
transform 1 0 1170 0 1 850
box 1170 850 1354 918
use cut_M1M4_2x1 
transform 1 0 1530 0 1 770
box 1530 770 1714 838
use cut_M1M4_2x1 
transform 1 0 1170 0 1 210
box 1170 210 1354 278
use cut_M1M4_2x1 
transform 1 0 1170 0 1 370
box 1170 370 1354 438
use cut_M1M4_2x1 
transform 1 0 1170 0 1 850
box 1170 850 1354 918
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1010
box 1170 1010 1354 1078
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1490
box 1170 1490 1354 1558
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1650
box 1170 1650 1354 1718
use cut_M1M4_2x1 
transform 1 0 1170 0 1 2130
box 1170 2130 1354 2198
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
<< labels >>
flabel locali s 1890 120 2070 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 630 1490 810 1550 0 FreeSans 400 0 0 0 N1
port 3 nsew
flabel locali s 630 1810 810 1870 0 FreeSans 400 0 0 0 N2
port 4 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 CI
port 5 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 CK
port 6 nsew
flabel locali s 630 2130 810 2190 0 FreeSans 400 0 0 0 CO
port 7 nsew
flabel locali s 270 2050 450 2110 0 FreeSans 400 0 0 0 VMR
port 8 nsew
flabel m3 s 1170 0 1354 2240 0 FreeSans 400 0 0 0 AVDD
port 9 nsew
flabel m3 s 630 0 814 2240 0 FreeSans 400 0 0 0 AVSS
port 10 nsew
<< end >>
