magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 10560
<< locali >>
rect 360 4610 498 4670
rect 498 4050 720 4110
rect 498 4050 558 4670
rect 360 5890 498 5950
rect 498 5330 720 5390
rect 498 5330 558 5950
rect 1422 3970 1620 4030
rect 1260 3730 1422 3790
rect 1422 3730 1482 4030
rect 360 8130 498 8190
rect 498 7890 720 7950
rect 498 7890 558 8190
rect 330 8130 390 8510
rect 390 9030 498 9090
rect 498 8850 720 8910
rect 498 8850 558 9090
rect 390 9090 450 9150
rect 390 9350 498 9410
rect 498 9170 720 9230
rect 498 9170 558 9410
rect 390 9410 450 9470
rect 360 10050 498 10110
rect 498 9650 720 9710
rect 498 9650 558 10110
rect 1260 5970 1398 6030
rect 1398 6530 1620 6590
rect 1398 5970 1458 6590
<< m1 >>
rect 360 5250 498 5310
rect 498 2770 720 2830
rect 498 2770 558 5318
rect 1620 7810 1758 7870
rect 1260 690 1758 750
rect 1758 690 1818 7878
rect 360 8770 498 8830
rect 498 7570 720 7630
rect 498 7570 558 8838
rect 1260 4690 1398 4750
rect 1398 7170 1620 7230
rect 1398 4690 1458 7238
<< m3 >>
rect 1712 4370 1772 6474
rect 1170 0 1354 10560
rect 630 0 814 10560
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use SARMRYX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 1980 3840
use SWX2_CV XA2
transform 1 0 0 0 1 3840
box 0 3840 1980 4480
use SWX2_CV XA3
transform 1 0 0 0 1 4480
box 0 4480 1980 5120
use SWX2_CV XA4
transform 1 0 0 0 1 5120
box 0 5120 1980 5760
use SWX2_CV XA5
transform 1 0 0 0 1 5760
box 0 5760 1980 6400
use SARCEX1_CV XA6
transform 1 0 0 0 1 6400
box 0 6400 1980 7680
use IVX1_CV XA7
transform 1 0 0 0 1 7680
box 0 7680 1980 8000
use IVX1_CV XA8
transform 1 0 0 0 1 8000
box 0 8000 1980 8320
use NDX1_CV XA9
transform 1 0 0 0 1 8320
box 0 8320 1980 8960
use IVX1_CV XA10
transform 1 0 0 0 1 8960
box 0 8960 1980 9280
use NRX1_CV XA11
transform 1 0 0 0 1 9280
box 0 9280 1980 9920
use IVX1_CV XA12
transform 1 0 0 0 1 9920
box 0 9920 1980 10240
use TAPCELLB_CV XA13
transform 1 0 0 0 1 10240
box 0 10240 1980 10560
use DMY_CV XA14
transform 1 0 0 0 1 10560
box 0 10560 0 10560
use cut_M1M2_2x1 
transform 1 0 270 0 1 5250
box 270 5250 454 5318
use cut_M1M2_2x1 
transform 1 0 630 0 1 2770
box 630 2770 814 2838
use cut_M1M2_2x1 
transform 1 0 1530 0 1 7810
box 1530 7810 1714 7878
use cut_M1M2_2x1 
transform 1 0 1170 0 1 690
box 1170 690 1354 758
use cut_M1M2_2x1 
transform 1 0 270 0 1 8770
box 270 8770 454 8838
use cut_M1M2_2x1 
transform 1 0 630 0 1 7570
box 630 7570 814 7638
use cut_M1M2_2x1 
transform 1 0 1170 0 1 4690
box 1170 4690 1354 4758
use cut_M1M2_2x1 
transform 1 0 1530 0 1 7170
box 1530 7170 1714 7238
use cut_M1M4_2x1 
transform 1 0 266 0 1 4606
box 266 4606 450 4674
use cut_M1M4_1x2 
transform 1 0 946 0 1 4628
box 946 4628 1014 4812
use cut_M1M4_1x2 
transform 1 0 1082 0 1 5268
box 1082 5268 1150 5452
use cut_M1M4_1x2 
transform 1 0 1218 0 1 5908
box 1218 5908 1286 6092
use cut_M2M3_2x1 
transform 1 0 1166 0 1 686
box 1166 686 1350 754
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
<< labels >>
flabel m2 s 266 2046 450 2114 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1530 3650 1710 3710 0 FreeSans 400 0 0 0 RST_N
port 2 nsew
flabel m2 s 266 446 450 514 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 270 3010 450 3070 0 FreeSans 400 0 0 0 CMP_ON
port 4 nsew
flabel m2 s 1166 686 1350 754 0 FreeSans 400 0 0 0 ENO
port 5 nsew
flabel m3 s 266 4606 450 4674 0 FreeSans 400 0 0 0 CN1
port 6 nsew
flabel m3 s 946 4628 1014 4812 0 FreeSans 400 0 0 0 CP1
port 7 nsew
flabel m3 s 1082 5268 1150 5452 0 FreeSans 400 0 0 0 CP0
port 8 nsew
flabel m3 s 1218 5908 1286 6092 0 FreeSans 400 0 0 0 CN0
port 9 nsew
flabel locali s 270 9730 450 9790 0 FreeSans 400 0 0 0 CEIN
port 10 nsew
flabel locali s 1170 10130 1350 10190 0 FreeSans 400 0 0 0 CEO
port 11 nsew
flabel locali s 270 6850 450 6910 0 FreeSans 400 0 0 0 CKS
port 12 nsew
flabel locali s 630 8210 810 8270 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 1650 4370 1834 4554 0 FreeSans 400 0 0 0 VREF
port 14 nsew
flabel m3 s 1170 0 1354 10560 0 FreeSans 400 0 0 0 AVDD
port 15 nsew
flabel m3 s 630 0 814 10560 0 FreeSans 400 0 0 0 AVSS
port 16 nsew
<< end >>
