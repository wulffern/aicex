magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 4104 2860
<< ppolyres >>
rect 162 -110 270 110
rect 378 -110 486 110
rect 594 -110 702 110
rect 810 -110 918 110
rect 1026 -110 1134 110
rect 1242 -110 1350 110
rect 1458 -110 1566 110
rect 1674 -110 1782 110
rect 1890 -110 1998 110
rect 2106 -110 2214 110
rect 2322 -110 2430 110
rect 2538 -110 2646 110
rect 2754 -110 2862 110
rect 2970 -110 3078 110
rect 3186 -110 3294 110
rect 3402 -110 3510 110
rect 3618 -110 3726 110
rect 3834 -110 3942 110
rect 162 110 270 330
rect 378 110 486 330
rect 594 110 702 330
rect 810 110 918 330
rect 1026 110 1134 330
rect 1242 110 1350 330
rect 1458 110 1566 330
rect 1674 110 1782 330
rect 1890 110 1998 330
rect 2106 110 2214 330
rect 2322 110 2430 330
rect 2538 110 2646 330
rect 2754 110 2862 330
rect 2970 110 3078 330
rect 3186 110 3294 330
rect 3402 110 3510 330
rect 3618 110 3726 330
rect 3834 110 3942 330
rect 162 330 270 550
rect 378 330 486 550
rect 594 330 702 550
rect 810 330 918 550
rect 1026 330 1134 550
rect 1242 330 1350 550
rect 1458 330 1566 550
rect 1674 330 1782 550
rect 1890 330 1998 550
rect 2106 330 2214 550
rect 2322 330 2430 550
rect 2538 330 2646 550
rect 2754 330 2862 550
rect 2970 330 3078 550
rect 3186 330 3294 550
rect 3402 330 3510 550
rect 3618 330 3726 550
rect 3834 330 3942 550
rect 162 550 270 770
rect 378 550 486 770
rect 594 550 702 770
rect 810 550 918 770
rect 1026 550 1134 770
rect 1242 550 1350 770
rect 1458 550 1566 770
rect 1674 550 1782 770
rect 1890 550 1998 770
rect 2106 550 2214 770
rect 2322 550 2430 770
rect 2538 550 2646 770
rect 2754 550 2862 770
rect 2970 550 3078 770
rect 3186 550 3294 770
rect 3402 550 3510 770
rect 3618 550 3726 770
rect 3834 550 3942 770
rect 162 770 270 990
rect 378 770 486 990
rect 594 770 702 990
rect 810 770 918 990
rect 1026 770 1134 990
rect 1242 770 1350 990
rect 1458 770 1566 990
rect 1674 770 1782 990
rect 1890 770 1998 990
rect 2106 770 2214 990
rect 2322 770 2430 990
rect 2538 770 2646 990
rect 2754 770 2862 990
rect 2970 770 3078 990
rect 3186 770 3294 990
rect 3402 770 3510 990
rect 3618 770 3726 990
rect 3834 770 3942 990
rect 162 990 270 1210
rect 378 990 486 1210
rect 594 990 702 1210
rect 810 990 918 1210
rect 1026 990 1134 1210
rect 1242 990 1350 1210
rect 1458 990 1566 1210
rect 1674 990 1782 1210
rect 1890 990 1998 1210
rect 2106 990 2214 1210
rect 2322 990 2430 1210
rect 2538 990 2646 1210
rect 2754 990 2862 1210
rect 2970 990 3078 1210
rect 3186 990 3294 1210
rect 3402 990 3510 1210
rect 3618 990 3726 1210
rect 3834 990 3942 1210
rect 162 1210 270 1430
rect 378 1210 486 1430
rect 594 1210 702 1430
rect 810 1210 918 1430
rect 1026 1210 1134 1430
rect 1242 1210 1350 1430
rect 1458 1210 1566 1430
rect 1674 1210 1782 1430
rect 1890 1210 1998 1430
rect 2106 1210 2214 1430
rect 2322 1210 2430 1430
rect 2538 1210 2646 1430
rect 2754 1210 2862 1430
rect 2970 1210 3078 1430
rect 3186 1210 3294 1430
rect 3402 1210 3510 1430
rect 3618 1210 3726 1430
rect 3834 1210 3942 1430
rect 162 1430 270 1650
rect 378 1430 486 1650
rect 594 1430 702 1650
rect 810 1430 918 1650
rect 1026 1430 1134 1650
rect 1242 1430 1350 1650
rect 1458 1430 1566 1650
rect 1674 1430 1782 1650
rect 1890 1430 1998 1650
rect 2106 1430 2214 1650
rect 2322 1430 2430 1650
rect 2538 1430 2646 1650
rect 2754 1430 2862 1650
rect 2970 1430 3078 1650
rect 3186 1430 3294 1650
rect 3402 1430 3510 1650
rect 3618 1430 3726 1650
rect 3834 1430 3942 1650
rect 162 1650 270 1870
rect 378 1650 486 1870
rect 594 1650 702 1870
rect 810 1650 918 1870
rect 1026 1650 1134 1870
rect 1242 1650 1350 1870
rect 1458 1650 1566 1870
rect 1674 1650 1782 1870
rect 1890 1650 1998 1870
rect 2106 1650 2214 1870
rect 2322 1650 2430 1870
rect 2538 1650 2646 1870
rect 2754 1650 2862 1870
rect 2970 1650 3078 1870
rect 3186 1650 3294 1870
rect 3402 1650 3510 1870
rect 3618 1650 3726 1870
rect 3834 1650 3942 1870
rect 162 1870 270 2090
rect 378 1870 486 2090
rect 594 1870 702 2090
rect 810 1870 918 2090
rect 1026 1870 1134 2090
rect 1242 1870 1350 2090
rect 1458 1870 1566 2090
rect 1674 1870 1782 2090
rect 1890 1870 1998 2090
rect 2106 1870 2214 2090
rect 2322 1870 2430 2090
rect 2538 1870 2646 2090
rect 2754 1870 2862 2090
rect 2970 1870 3078 2090
rect 3186 1870 3294 2090
rect 3402 1870 3510 2090
rect 3618 1870 3726 2090
rect 3834 1870 3942 2090
rect 162 2090 270 2310
rect 378 2090 486 2310
rect 594 2090 702 2310
rect 810 2090 918 2310
rect 1026 2090 1134 2310
rect 1242 2090 1350 2310
rect 1458 2090 1566 2310
rect 1674 2090 1782 2310
rect 1890 2090 1998 2310
rect 2106 2090 2214 2310
rect 2322 2090 2430 2310
rect 2538 2090 2646 2310
rect 2754 2090 2862 2310
rect 2970 2090 3078 2310
rect 3186 2090 3294 2310
rect 3402 2090 3510 2310
rect 3618 2090 3726 2310
rect 3834 2090 3942 2310
rect 162 2310 270 2530
rect 378 2310 486 2530
rect 594 2310 702 2530
rect 810 2310 918 2530
rect 1026 2310 1134 2530
rect 1242 2310 1350 2530
rect 1458 2310 1566 2530
rect 1674 2310 1782 2530
rect 1890 2310 1998 2530
rect 2106 2310 2214 2530
rect 2322 2310 2430 2530
rect 2538 2310 2646 2530
rect 2754 2310 2862 2530
rect 2970 2310 3078 2530
rect 3186 2310 3294 2530
rect 3402 2310 3510 2530
rect 3618 2310 3726 2530
rect 3834 2310 3942 2530
<< poly >>
rect -54 -110 54 110
rect 4050 -110 4158 110
rect -54 110 54 330
rect 4050 110 4158 330
rect -54 330 54 550
rect 4050 330 4158 550
rect -54 550 54 770
rect 4050 550 4158 770
rect -54 770 54 990
rect 4050 770 4158 990
rect -54 990 54 1210
rect 4050 990 4158 1210
rect -54 1210 54 1430
rect 4050 1210 4158 1430
rect -54 1430 54 1650
rect 4050 1430 4158 1650
rect -54 1650 54 1870
rect 4050 1650 4158 1870
rect -54 1870 54 2090
rect 4050 1870 4158 2090
rect -54 2090 54 2310
rect 4050 2090 4158 2310
rect -54 2310 54 2530
rect 4050 2310 4158 2530
<< xpolycontact >>
rect 162 -110 270 110
rect 378 -110 486 110
rect 594 -110 702 110
rect 810 -110 918 110
rect 1026 -110 1134 110
rect 1242 -110 1350 110
rect 1458 -110 1566 110
rect 1674 -110 1782 110
rect 1890 -110 1998 110
rect 2106 -110 2214 110
rect 2322 -110 2430 110
rect 2538 -110 2646 110
rect 2754 -110 2862 110
rect 2970 -110 3078 110
rect 3186 -110 3294 110
rect 3402 -110 3510 110
rect 3618 -110 3726 110
rect 3834 -110 3942 110
rect 162 110 270 330
rect 378 110 486 330
rect 594 110 702 330
rect 810 110 918 330
rect 1026 110 1134 330
rect 1242 110 1350 330
rect 1458 110 1566 330
rect 1674 110 1782 330
rect 1890 110 1998 330
rect 2106 110 2214 330
rect 2322 110 2430 330
rect 2538 110 2646 330
rect 2754 110 2862 330
rect 2970 110 3078 330
rect 3186 110 3294 330
rect 3402 110 3510 330
rect 3618 110 3726 330
rect 3834 110 3942 330
rect 162 2090 270 2310
rect 378 2090 486 2310
rect 594 2090 702 2310
rect 810 2090 918 2310
rect 1026 2090 1134 2310
rect 1242 2090 1350 2310
rect 1458 2090 1566 2310
rect 1674 2090 1782 2310
rect 1890 2090 1998 2310
rect 2106 2090 2214 2310
rect 2322 2090 2430 2310
rect 2538 2090 2646 2310
rect 2754 2090 2862 2310
rect 2970 2090 3078 2310
rect 3186 2090 3294 2310
rect 3402 2090 3510 2310
rect 3618 2090 3726 2310
rect 3834 2090 3942 2310
rect 162 2310 270 2530
rect 378 2310 486 2530
rect 594 2310 702 2530
rect 810 2310 918 2530
rect 1026 2310 1134 2530
rect 1242 2310 1350 2530
rect 1458 2310 1566 2530
rect 1674 2310 1782 2530
rect 1890 2310 1998 2530
rect 2106 2310 2214 2530
rect 2322 2310 2430 2530
rect 2538 2310 2646 2530
rect 2754 2310 2862 2530
rect 2970 2310 3078 2530
rect 3186 2310 3294 2530
rect 3402 2310 3510 2530
rect 3618 2310 3726 2530
rect 3834 2310 3942 2530
<< locali >>
rect 162 -110 486 110
rect 594 -110 918 110
rect 1026 -110 1350 110
rect 1458 -110 1782 110
rect 1890 -110 2214 110
rect 2322 -110 2646 110
rect 2754 -110 3078 110
rect 3186 -110 3510 110
rect 3618 -110 3942 110
rect 162 110 486 330
rect 594 110 918 330
rect 1026 110 1350 330
rect 1458 110 1782 330
rect 1890 110 2214 330
rect 2322 110 2646 330
rect 2754 110 3078 330
rect 3186 110 3510 330
rect 3618 110 3942 330
rect 162 2090 270 2310
rect 378 2090 486 2310
rect 594 2090 702 2310
rect 810 2090 918 2310
rect 1026 2090 1134 2310
rect 1242 2090 1350 2310
rect 1458 2090 1566 2310
rect 1674 2090 1782 2310
rect 1890 2090 1998 2310
rect 2106 2090 2214 2310
rect 2322 2090 2430 2310
rect 2538 2090 2646 2310
rect 2754 2090 2862 2310
rect 2970 2090 3078 2310
rect 3186 2090 3294 2310
rect 3402 2090 3510 2310
rect 3618 2090 3726 2310
rect 3834 2090 3942 2310
rect 162 2310 270 2530
rect 378 2310 486 2530
rect 594 2310 702 2530
rect 810 2310 918 2530
rect 1026 2310 1134 2530
rect 1242 2310 1350 2530
rect 1458 2310 1566 2530
rect 1674 2310 1782 2530
rect 1890 2310 1998 2530
rect 2106 2310 2214 2530
rect 2322 2310 2430 2530
rect 2538 2310 2646 2530
rect 2754 2310 2862 2530
rect 2970 2310 3078 2530
rect 3186 2310 3294 2530
rect 3402 2310 3510 2530
rect 3618 2310 3726 2530
rect 3834 2310 3942 2530
rect 162 2530 270 2750
rect 378 2530 486 2750
rect 594 2530 702 2750
rect 810 2530 918 2750
rect 1026 2530 1134 2750
rect 1242 2530 1350 2750
rect 1458 2530 1566 2750
rect 1674 2530 1782 2750
rect 1890 2530 1998 2750
rect 2106 2530 2214 2750
rect 2322 2530 2430 2750
rect 2538 2530 2646 2750
rect 2754 2530 2862 2750
rect 2970 2530 3078 2750
rect 3186 2530 3294 2750
rect 3402 2530 3510 2750
rect 3618 2530 3726 2750
rect 3834 2530 3942 2750
rect -54 2750 270 2970
rect -54 2750 270 2970
rect 378 2750 702 2970
rect 810 2750 1134 2970
rect 1242 2750 1566 2970
rect 1674 2750 1998 2970
rect 2106 2750 2430 2970
rect 2538 2750 2862 2970
rect 2970 2750 3294 2970
rect 3402 2750 3726 2970
rect 3834 2750 4158 2970
rect 3834 2750 4158 2970
<< pwell >>
rect -54 -110 4158 2970
<< labels >>
flabel locali s -54 2750 270 2970 0 FreeSans 400 0 0 0 N
port 1 nsew
flabel locali s 3834 2750 4158 2970 0 FreeSans 400 0 0 0 P
port 2 nsew
<< end >>
