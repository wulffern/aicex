magic
tech sky130A
magscale 1 2
timestamp 1664582400
<< checkpaint >>
rect 0 0 3536 4236
<< locali >>
rect 16 16 3520 128
rect 16 16 3520 128
rect 16 16 128 4220
rect 16 4108 3520 4220
rect 3408 16 3520 4220
rect 16 16 3520 128
rect 2344 3438 2920 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 48 32 128 112
rect 128 32 208 112
rect 208 32 288 112
rect 288 32 368 112
rect 368 32 448 112
rect 448 32 528 112
rect 528 32 608 112
rect 608 32 688 112
rect 688 32 768 112
rect 768 32 848 112
rect 848 32 928 112
rect 928 32 1008 112
rect 1008 32 1088 112
rect 1088 32 1168 112
rect 1168 32 1248 112
rect 1248 32 1328 112
rect 1328 32 1408 112
rect 1408 32 1488 112
rect 1488 32 1568 112
rect 1568 32 1648 112
rect 1648 32 1728 112
rect 1728 32 1808 112
rect 1808 32 1888 112
rect 1888 32 1968 112
rect 1968 32 2048 112
rect 2048 32 2128 112
rect 2128 32 2208 112
rect 2208 32 2288 112
rect 2288 32 2368 112
rect 2368 32 2448 112
rect 2448 32 2528 112
rect 2528 32 2608 112
rect 2608 32 2688 112
rect 2688 32 2768 112
rect 2768 32 2848 112
rect 2848 32 2928 112
rect 2928 32 3008 112
rect 3008 32 3088 112
rect 3088 32 3168 112
rect 3168 32 3248 112
rect 3248 32 3328 112
rect 3328 32 3408 112
rect 3408 32 3488 112
rect 32 38 112 118
rect 32 118 112 198
rect 32 198 112 278
rect 32 278 112 358
rect 32 358 112 438
rect 32 438 112 518
rect 32 518 112 598
rect 32 598 112 678
rect 32 678 112 758
rect 32 758 112 838
rect 32 838 112 918
rect 32 918 112 998
rect 32 998 112 1078
rect 32 1078 112 1158
rect 32 1158 112 1238
rect 32 1238 112 1318
rect 32 1318 112 1398
rect 32 1398 112 1478
rect 32 1478 112 1558
rect 32 1558 112 1638
rect 32 1638 112 1718
rect 32 1718 112 1798
rect 32 1798 112 1878
rect 32 1878 112 1958
rect 32 1958 112 2038
rect 32 2038 112 2118
rect 32 2118 112 2198
rect 32 2198 112 2278
rect 32 2278 112 2358
rect 32 2358 112 2438
rect 32 2438 112 2518
rect 32 2518 112 2598
rect 32 2598 112 2678
rect 32 2678 112 2758
rect 32 2758 112 2838
rect 32 2838 112 2918
rect 32 2918 112 2998
rect 32 2998 112 3078
rect 32 3078 112 3158
rect 32 3158 112 3238
rect 32 3238 112 3318
rect 32 3318 112 3398
rect 32 3398 112 3478
rect 32 3478 112 3558
rect 32 3558 112 3638
rect 32 3638 112 3718
rect 32 3718 112 3798
rect 32 3798 112 3878
rect 32 3878 112 3958
rect 32 3958 112 4038
rect 32 4038 112 4118
rect 32 4118 112 4198
rect 48 4124 128 4204
rect 128 4124 208 4204
rect 208 4124 288 4204
rect 288 4124 368 4204
rect 368 4124 448 4204
rect 448 4124 528 4204
rect 528 4124 608 4204
rect 608 4124 688 4204
rect 688 4124 768 4204
rect 768 4124 848 4204
rect 848 4124 928 4204
rect 928 4124 1008 4204
rect 1008 4124 1088 4204
rect 1088 4124 1168 4204
rect 1168 4124 1248 4204
rect 1248 4124 1328 4204
rect 1328 4124 1408 4204
rect 1408 4124 1488 4204
rect 1488 4124 1568 4204
rect 1568 4124 1648 4204
rect 1648 4124 1728 4204
rect 1728 4124 1808 4204
rect 1808 4124 1888 4204
rect 1888 4124 1968 4204
rect 1968 4124 2048 4204
rect 2048 4124 2128 4204
rect 2128 4124 2208 4204
rect 2208 4124 2288 4204
rect 2288 4124 2368 4204
rect 2368 4124 2448 4204
rect 2448 4124 2528 4204
rect 2528 4124 2608 4204
rect 2608 4124 2688 4204
rect 2688 4124 2768 4204
rect 2768 4124 2848 4204
rect 2848 4124 2928 4204
rect 2928 4124 3008 4204
rect 3008 4124 3088 4204
rect 3088 4124 3168 4204
rect 3168 4124 3248 4204
rect 3248 4124 3328 4204
rect 3328 4124 3408 4204
rect 3408 4124 3488 4204
rect 3424 38 3504 118
rect 3424 118 3504 198
rect 3424 198 3504 278
rect 3424 278 3504 358
rect 3424 358 3504 438
rect 3424 438 3504 518
rect 3424 518 3504 598
rect 3424 598 3504 678
rect 3424 678 3504 758
rect 3424 758 3504 838
rect 3424 838 3504 918
rect 3424 918 3504 998
rect 3424 998 3504 1078
rect 3424 1078 3504 1158
rect 3424 1158 3504 1238
rect 3424 1238 3504 1318
rect 3424 1318 3504 1398
rect 3424 1398 3504 1478
rect 3424 1478 3504 1558
rect 3424 1558 3504 1638
rect 3424 1638 3504 1718
rect 3424 1718 3504 1798
rect 3424 1798 3504 1878
rect 3424 1878 3504 1958
rect 3424 1958 3504 2038
rect 3424 2038 3504 2118
rect 3424 2118 3504 2198
rect 3424 2198 3504 2278
rect 3424 2278 3504 2358
rect 3424 2358 3504 2438
rect 3424 2438 3504 2518
rect 3424 2518 3504 2598
rect 3424 2598 3504 2678
rect 3424 2678 3504 2758
rect 3424 2758 3504 2838
rect 3424 2838 3504 2918
rect 3424 2918 3504 2998
rect 3424 2998 3504 3078
rect 3424 3078 3504 3158
rect 3424 3158 3504 3238
rect 3424 3238 3504 3318
rect 3424 3318 3504 3398
rect 3424 3398 3504 3478
rect 3424 3478 3504 3558
rect 3424 3558 3504 3638
rect 3424 3638 3504 3718
rect 3424 3718 3504 3798
rect 3424 3798 3504 3878
rect 3424 3878 3504 3958
rect 3424 3958 3504 4038
rect 3424 4038 3504 4118
rect 3424 4118 3504 4198
<< ptap >>
rect 0 0 3536 144
rect 0 0 144 4236
rect 0 4092 3536 4236
rect 3392 0 3536 4236
use SUNTR_RES4 XA1
transform 1 0 688 0 1 688
box 688 688 2848 3548
<< labels >>
flabel locali s 16 16 3520 128 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 2344 3438 2920 3658 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
