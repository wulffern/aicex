
.lib Rt

*.include "../../../models/skywater-pdk-libs-sky130_fd_pr/models/r+c/res_typical__cap_typical.spice"
*.include "../../../models/skywater-pdk-libs-sky130_fd_pr/models/r+c/res_typical__cap_typical__lin.spice"

*.include "../../../models/skywater-pdk-libs-sky130_fd_pr/cells/res_xhigh_po/sky130_fd_pr__res_xhigh_po.model.spice"
*.include "../../../models/skywater-pdk-libs-sky130_fd_pr/cells/res_high_po/sky130_fd_pr__res_high_po.model.spice"



.endl

.lib Rl

* TODO does not seem like there is a high res corner



.endl

.lib Rh

* TODO does not seem like there is a high res corner



.endl
