magic
tech sky130A
magscale 1 2
timestamp 1664582400
<< checkpaint >>
rect 0 0 1260 528
<< ndiff >>
rect 756 132 972 220
rect 756 220 972 308
rect 756 308 972 396
<< ptap >>
rect -108 -44 108 44
rect -108 44 108 132
rect -108 132 108 220
rect -108 220 108 308
rect -108 308 108 396
rect -108 396 108 484
rect -108 484 108 572
<< poly >>
rect 324 -36 1044 36
rect 324 228 1044 300
rect 324 492 1044 564
rect 324 220 540 308
<< locali >>
rect 324 234 540 294
rect -108 -44 108 44
rect -108 44 108 132
rect -108 132 108 220
rect 756 146 972 206
rect 756 146 972 206
rect -108 220 108 308
rect -108 220 108 308
rect 324 234 540 294
rect -108 308 108 396
rect 756 322 972 382
rect 756 322 972 382
rect -108 396 108 484
rect -108 484 108 572
<< pcontact >>
rect 348 242 396 264
rect 348 264 396 286
rect 396 242 468 264
rect 396 264 468 286
rect 468 242 516 264
rect 468 264 516 286
<< ptapc >>
rect -36 132 36 220
rect -36 308 36 396
<< ndcontact >>
rect 780 154 828 176
rect 780 176 828 198
rect 828 154 900 176
rect 828 176 900 198
rect 900 154 948 176
rect 900 176 948 198
rect 780 330 828 352
rect 780 352 828 374
rect 828 330 900 352
rect 828 352 900 374
rect 900 330 948 352
rect 900 352 948 374
<< pwell >>
rect -180 -132 1260 660
<< labels >>
flabel locali s 324 234 540 294 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 756 146 972 206 0 FreeSans 400 0 0 0 S
port 3 nsew
flabel locali s -108 220 108 308 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 756 322 972 382 0 FreeSans 400 0 0 0 D
port 1 nsew
<< end >>
