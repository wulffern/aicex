

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../lib/SUN_TR_SKY130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------

VSS VSS 0 dc 0
INN 0 N1 dc 1.0u

XM1 N1 N1 VSS VSS NCH

.probe v(n1)

.control
set color0=white
set color1=black
unset askquit
*set filetype=ascii
*set appendwrite=1
dc inn 0.01u 100u 0.01u

write

quit
.endc
.end
