magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 14712 11040
<< locali >>
rect 14088 384 14328 10656
rect 384 384 14328 624
rect 384 10416 14328 10656
rect 384 384 624 10656
rect 14088 384 14328 10656
rect 14472 0 14712 11040
rect 0 0 14712 240
rect 0 10800 14712 11040
rect 0 0 240 11040
rect 14472 0 14712 11040
rect 1632 2410 1800 2470
rect 1632 2586 1800 2646
rect 1632 3114 1800 3174
rect 1800 2410 1860 3174
rect 3252 826 3420 886
rect 3252 2058 3420 2118
rect 3252 3290 3420 3350
rect 3252 4522 3420 4582
rect 3252 5754 3420 5814
rect 3420 826 3480 5814
<< m1 >>
rect 1524 384 1740 886
rect 660 384 876 988
rect 660 384 876 2748
rect 660 384 876 3276
rect 3144 0 3360 886
rect 2280 0 2496 988
rect 2820 5842 2988 5902
rect 2988 1002 3252 1062
rect 2820 3378 2988 3438
rect 2820 4610 2988 4670
rect 1632 3290 2988 3350
rect 2988 1002 3048 5902
<< m3 >>
rect 8796 384 9012 812
rect 3252 3466 3432 3542
rect 3252 4698 3432 4774
rect 3252 5930 3432 6006
rect 3432 1604 8904 1680
rect 3432 2660 8904 2736
rect 3432 3716 8904 3792
rect 3432 4772 8904 4848
rect 3432 5828 8904 5904
rect 3432 6884 8904 6960
rect 3432 7940 8904 8016
rect 3432 8996 8904 9072
rect 3432 10052 8904 10128
rect 3432 1604 3508 10128
rect 8904 724 14196 800
rect 8904 1780 14196 1856
rect 8904 2836 14196 2912
rect 8904 3892 14196 3968
rect 8904 4948 14196 5024
rect 8904 6004 14196 6080
rect 8904 7060 14196 7136
rect 8904 8116 14196 8192
rect 8904 9172 14196 9248
rect 14196 724 14272 9248
<< m2 >>
rect 2820 914 2992 990
rect 1632 2762 2992 2838
rect 2992 2234 3252 2310
rect 2820 2146 2992 2222
rect 2992 914 3068 2838
rect 0 2674 216 2734
rect 0 3202 216 3262
rect 0 3466 216 3526
rect 0 914 216 974
rect 0 914 216 974
rect 952 914 1200 990
rect 108 914 952 990
rect 952 914 1028 990
rect 0 2674 216 2734
rect 952 2674 1200 2750
rect 108 2674 952 2750
rect 952 2674 1028 2750
rect 0 3202 216 3262
rect 952 3202 1200 3278
rect 108 3202 952 3278
rect 952 3202 1028 3278
rect 0 3466 216 3526
rect 3004 3466 3252 3542
rect 108 3466 3004 3542
rect 3004 3466 3080 3542
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa10
transform 1 0 768 0 1 768
box 768 768 2028 2528
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa20
transform 1 0 768 0 1 2528
box 768 2528 2028 3056
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa40
transform 1 0 768 0 1 3056
box 768 3056 2028 3584
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc10
transform -1 0 3648 0 1 768
box 3648 768 4908 2000
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc20
transform -1 0 3648 0 1 2000
box 3648 2000 4908 3232
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_00
transform -1 0 3648 0 1 3232
box 3648 3232 4908 4464
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_10
transform -1 0 3648 0 1 4464
box 3648 4464 4908 5696
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_20
transform -1 0 3648 0 1 5696
box 3648 5696 4908 6928
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd20
transform 1 0 3792 0 1 768
box 3792 768 13944 1824
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd30
transform 1 0 3792 0 1 1824
box 3792 1824 13944 2880
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd31
transform 1 0 3792 0 1 2880
box 3792 2880 13944 3936
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd32
transform 1 0 3792 0 1 3936
box 3792 3936 13944 4992
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd33
transform 1 0 3792 0 1 4992
box 3792 4992 13944 6048
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd34
transform 1 0 3792 0 1 6048
box 3792 6048 13944 7104
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd35
transform 1 0 3792 0 1 7104
box 3792 7104 13944 8160
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd36
transform 1 0 3792 0 1 8160
box 3792 8160 13944 9216
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd37
transform 1 0 3792 0 1 9216
box 3792 9216 13944 10272
use cut_M1M2_2x1 
transform 1 0 1540 0 1 826
box 1540 826 1724 894
use cut_M1M2_2x1 
transform 1 0 1540 0 1 384
box 1540 384 1724 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 900
box 676 900 860 968
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 2660
box 676 2660 860 2728
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 3188
box 676 3188 860 3256
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M4_2x1 
transform 1 0 8804 0 1 384
box 8804 384 9004 460
use cut_M1M2_2x1 
transform 1 0 3160 0 1 826
box 3160 826 3344 894
use cut_M1M2_2x1 
transform 1 0 3160 0 1 0
box 3160 0 3344 68
use cut_M1M2_2x1 
transform 1 0 2296 0 1 900
box 2296 900 2480 968
use cut_M1M2_2x1 
transform 1 0 2296 0 1 0
box 2296 0 2480 68
use cut_M1M2_2x1 
transform 1 0 2712 0 1 5842
box 2712 5842 2896 5910
use cut_M1M2_2x1 
transform 1 0 3144 0 1 1002
box 3144 1002 3328 1070
use cut_M1M2_2x1 
transform 1 0 2712 0 1 3378
box 2712 3378 2896 3446
use cut_M1M2_2x1 
transform 1 0 2712 0 1 4610
box 2712 4610 2896 4678
use cut_M1M2_2x1 
transform 1 0 1524 0 1 3290
box 1524 3290 1708 3358
use cut_M1M3_2x1 
transform 1 0 2712 0 1 914
box 2712 914 2912 990
use cut_M1M3_2x1 
transform 1 0 1524 0 1 2762
box 1524 2762 1724 2838
use cut_M1M3_2x1 
transform 1 0 3144 0 1 2234
box 3144 2234 3344 2310
use cut_M1M3_2x1 
transform 1 0 2712 0 1 2146
box 2712 2146 2912 2222
use cut_M1M4_2x1 
transform 1 0 3144 0 1 3466
box 3144 3466 3344 3542
use cut_M1M4_2x1 
transform 1 0 3144 0 1 4698
box 3144 4698 3344 4774
use cut_M1M4_2x1 
transform 1 0 3144 0 1 5930
box 3144 5930 3344 6006
use cut_M1M3_2x1 
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M3_2x1 
transform 1 0 1108 0 1 2674
box 1108 2674 1308 2750
use cut_M1M3_2x1 
transform 1 0 1108 0 1 3202
box 1108 3202 1308 3278
use cut_M1M3_2x1 
transform 1 0 3160 0 1 3466
box 3160 3466 3360 3542
<< labels >>
flabel locali s 14088 384 14328 10656 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 14472 0 14712 11040 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 0 2674 216 2734 0 FreeSans 400 0 0 0 VFB
port 2 nsew
flabel m2 s 0 3202 216 3262 0 FreeSans 400 0 0 0 VI
port 3 nsew
flabel m2 s 0 3466 216 3526 0 FreeSans 400 0 0 0 VO
port 4 nsew
flabel m2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew
<< end >>
