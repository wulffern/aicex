magic
tech sky130A
magscale 1 2
timestamp 1658775803
<< checkpaint >>
rect -2284 0 26372 55382
<< m3 >>
rect 9100 33880 26178 33956
rect 9100 34268 26178 34344
rect 24104 34648 24180 42152
rect 24384 34648 24460 49896
rect 3944 34732 4020 45664
rect 4824 34926 4900 45664
rect 8984 35120 9060 45664
rect -216 35314 -140 45664
rect -216 35314 -140 45664
rect 13432 35508 13508 45690
rect 13432 35508 13508 45690
rect 18472 35702 18548 45690
rect 18472 35702 18548 45690
rect 10579 35896 10655 45690
rect 10579 35896 10655 45690
rect 15619 36090 15695 45690
rect 15619 36090 15695 45690
rect 499 36284 575 45690
rect 5539 36478 5615 45690
rect 5539 36478 5615 45690
rect 3352 36672 3428 45690
rect 3352 36672 3428 45690
rect 8392 36866 8468 45690
rect 8392 36866 8468 45690
rect 659 37060 735 47098
rect 8232 37254 8308 47098
rect 5699 37448 5775 47098
rect 3192 37642 3268 47098
rect 10914 37836 10990 48506
rect 13098 38030 13174 48506
rect 15954 38224 16030 48506
rect 8058 38418 8134 48506
rect 3018 38612 3094 48506
rect 834 38806 910 48506
rect 18138 39000 18214 48506
rect 5874 39194 5950 48506
rect 11072 50 11272 126
rect 12816 50 13016 126
rect 20659 45690 20735 45890
rect 1568 44704 1768 44904
rect 8856 0 9056 5280
rect 9648 0 9848 5280
<< m2 >>
rect 14872 33374 14948 33956
rect 9100 33374 9176 34344
rect 3944 34656 14020 34732
rect 4824 34850 13660 34926
rect 8984 35044 13300 35120
rect -216 35238 14380 35314
rect 11304 35432 13508 35508
rect 11664 35626 18548 35702
rect 10579 35820 11200 35896
rect 11484 36014 15695 36090
rect 499 36208 9760 36284
rect 5539 36402 10480 36478
rect 3352 36596 10120 36672
rect 8392 36790 10840 36866
rect 659 36984 9940 37060
rect 8232 37178 11020 37254
rect 5699 37372 10660 37448
rect 3192 37566 10300 37642
rect 10914 37760 12940 37836
rect 12684 37954 13174 38030
rect 12504 38148 16030 38224
rect 8058 38342 13120 38418
rect 3018 38536 13840 38612
rect 834 38730 14200 38806
rect 12324 38924 18214 39000
rect 5874 39118 13480 39194
rect -216 40384 -16 40460
<< m4 >>
rect 24104 34268 24180 34648
rect 24384 33880 24460 34648
<< m1 >>
rect 13944 33314 14020 34656
rect 13584 33314 13660 34850
rect 13224 33314 13300 35044
rect 14304 33314 14380 35238
rect 11304 33314 11380 35432
rect 11664 33314 11740 35626
rect 11124 33314 11200 35820
rect 11484 33314 11560 36014
rect 9684 33314 9760 36208
rect 10404 33314 10480 36402
rect 10044 33314 10120 36596
rect 10764 33314 10840 36790
rect 9864 33314 9940 36984
rect 10944 33314 11020 37178
rect 10584 33314 10660 37372
rect 10224 33314 10300 37566
rect 12864 33314 12940 37760
rect 12684 33314 12760 37954
rect 12504 33314 12580 38148
rect 13044 33314 13120 38342
rect 13764 33314 13840 38536
rect 14124 33314 14200 38730
rect 12324 33314 12400 38924
rect 13404 33314 13480 39118
<< locali >>
rect 11072 2698 11288 2758
rect 11072 1290 11288 1350
rect 20360 51744 20576 51804
rect -232 50248 -16 50308
rect 10064 498 10280 558
use SARBSSW_CV XB1
transform -1 0 12044 0 1 0
box 12044 0 26372 5280
use SARBSSW_CV XB2
transform 1 0 12044 0 1 0
box 12044 0 26372 5280
use CDAC8_CV XDAC1
transform -1 0 11844 0 1 5474
box 11844 5474 23576 33374
use CDAC8_CV XDAC2
transform 1 0 12204 0 1 5474
box 12204 5474 23936 33374
use SARDIGEX4_CV XA0
transform 1 0 -556 0 1 39894
box -556 39894 1964 54326
use SARDIGEX4_CV XA1
transform -1 0 4484 0 1 39894
box 4484 39894 7004 54326
use SARDIGEX4_CV XA2
transform 1 0 4484 0 1 39894
box 4484 39894 7004 54326
use SARDIGEX4_CV XA3
transform -1 0 9524 0 1 39894
box 9524 39894 12044 54326
use SARDIGEX4_CV XA4
transform 1 0 9524 0 1 39894
box 9524 39894 12044 54326
use SARDIGEX4_CV XA5
transform -1 0 14564 0 1 39894
box 14564 39894 17084 54326
use SARDIGEX4_CV XA6
transform 1 0 14564 0 1 39894
box 14564 39894 17084 54326
use SARDIGEX4_CV XA7
transform -1 0 19604 0 1 39894
box 19604 39894 22124 54326
use SARDIGEX4_CV XA8
transform 1 0 19604 0 1 39894
box 19604 39894 22124 54326
use SARCMPX1_CV XA20
transform -1 0 24644 0 1 39894
box 24644 39894 27164 55382
use cut_M3M4_1x2 
transform 1 0 14872 0 1 33374
box 14872 33374 14948 33574
use cut_M3M4_2x1 
transform 1 0 14872 0 1 33880
box 14872 33880 15072 33956
use cut_M3M4_1x2 
transform 1 0 9100 0 1 33374
box 9100 33374 9176 33574
use cut_M3M4_2x1 
transform 1 0 9100 0 1 34268
box 9100 34268 9300 34344
use cut_M2M4_2x1 
transform 1 0 24104 0 1 42152
box 24104 42152 24304 42228
use cut_M4M5_2x1 
transform 1 0 24104 0 1 34268
box 24104 34268 24304 34344
use cut_M4M5_1x2 
transform 1 0 24104 0 1 34648
box 24104 34648 24180 34848
use cut_M3M4_2x1 
transform 1 0 24260 0 1 49896
box 24260 49896 24460 49972
use cut_M2M3_2x1 
transform 1 0 24104 0 1 49896
box 24104 49896 24304 49972
use cut_M4M5_2x1 
transform 1 0 24384 0 1 33880
box 24384 33880 24584 33956
use cut_M4M5_1x2 
transform 1 0 24384 0 1 34648
box 24384 34648 24460 34848
use cut_M3M4_1x2 
transform 1 0 3944 0 1 34594
box 3944 34594 4020 34794
use cut_M2M3_1x2 
transform 1 0 13936 0 1 34594
box 13936 34594 14012 34794
use cut_M3M4_1x2 
transform 1 0 4824 0 1 34788
box 4824 34788 4900 34988
use cut_M2M3_1x2 
transform 1 0 13576 0 1 34788
box 13576 34788 13652 34988
use cut_M3M4_1x2 
transform 1 0 8984 0 1 34982
box 8984 34982 9060 35182
use cut_M2M3_1x2 
transform 1 0 13216 0 1 34982
box 13216 34982 13292 35182
use cut_M3M4_1x2 
transform 1 0 -216 0 1 35176
box -216 35176 -140 35376
use cut_M2M3_1x2 
transform 1 0 14296 0 1 35176
box 14296 35176 14372 35376
use cut_M3M4_1x2 
transform 1 0 13432 0 1 35370
box 13432 35370 13508 35570
use cut_M2M3_1x2 
transform 1 0 11296 0 1 35370
box 11296 35370 11372 35570
use cut_M3M4_1x2 
transform 1 0 18472 0 1 35564
box 18472 35564 18548 35764
use cut_M2M3_1x2 
transform 1 0 11656 0 1 35564
box 11656 35564 11732 35764
use cut_M3M4_1x2 
transform 1 0 10579 0 1 35758
box 10579 35758 10655 35958
use cut_M2M3_1x2 
transform 1 0 11116 0 1 35758
box 11116 35758 11192 35958
use cut_M3M4_1x2 
transform 1 0 15619 0 1 35952
box 15619 35952 15695 36152
use cut_M2M3_1x2 
transform 1 0 11476 0 1 35952
box 11476 35952 11552 36152
use cut_M3M4_1x2 
transform 1 0 499 0 1 36146
box 499 36146 575 36346
use cut_M2M3_1x2 
transform 1 0 9676 0 1 36146
box 9676 36146 9752 36346
use cut_M3M4_1x2 
transform 1 0 5539 0 1 36340
box 5539 36340 5615 36540
use cut_M2M3_1x2 
transform 1 0 10396 0 1 36340
box 10396 36340 10472 36540
use cut_M3M4_1x2 
transform 1 0 3352 0 1 36534
box 3352 36534 3428 36734
use cut_M2M3_1x2 
transform 1 0 10036 0 1 36534
box 10036 36534 10112 36734
use cut_M3M4_1x2 
transform 1 0 8392 0 1 36728
box 8392 36728 8468 36928
use cut_M2M3_1x2 
transform 1 0 10756 0 1 36728
box 10756 36728 10832 36928
use cut_M3M4_1x2 
transform 1 0 659 0 1 36922
box 659 36922 735 37122
use cut_M2M3_1x2 
transform 1 0 9856 0 1 36922
box 9856 36922 9932 37122
use cut_M3M4_1x2 
transform 1 0 8232 0 1 37116
box 8232 37116 8308 37316
use cut_M2M3_1x2 
transform 1 0 10936 0 1 37116
box 10936 37116 11012 37316
use cut_M3M4_1x2 
transform 1 0 5699 0 1 37310
box 5699 37310 5775 37510
use cut_M2M3_1x2 
transform 1 0 10576 0 1 37310
box 10576 37310 10652 37510
use cut_M3M4_1x2 
transform 1 0 3192 0 1 37504
box 3192 37504 3268 37704
use cut_M2M3_1x2 
transform 1 0 10216 0 1 37504
box 10216 37504 10292 37704
use cut_M3M4_1x2 
transform 1 0 10914 0 1 37698
box 10914 37698 10990 37898
use cut_M2M3_1x2 
transform 1 0 12856 0 1 37698
box 12856 37698 12932 37898
use cut_M3M4_1x2 
transform 1 0 13098 0 1 37892
box 13098 37892 13174 38092
use cut_M2M3_1x2 
transform 1 0 12676 0 1 37892
box 12676 37892 12752 38092
use cut_M3M4_1x2 
transform 1 0 15954 0 1 38086
box 15954 38086 16030 38286
use cut_M2M3_1x2 
transform 1 0 12496 0 1 38086
box 12496 38086 12572 38286
use cut_M3M4_1x2 
transform 1 0 8058 0 1 38280
box 8058 38280 8134 38480
use cut_M2M3_1x2 
transform 1 0 13036 0 1 38280
box 13036 38280 13112 38480
use cut_M3M4_1x2 
transform 1 0 3018 0 1 38474
box 3018 38474 3094 38674
use cut_M2M3_1x2 
transform 1 0 13756 0 1 38474
box 13756 38474 13832 38674
use cut_M3M4_1x2 
transform 1 0 834 0 1 38668
box 834 38668 910 38868
use cut_M2M3_1x2 
transform 1 0 14116 0 1 38668
box 14116 38668 14192 38868
use cut_M3M4_1x2 
transform 1 0 18138 0 1 38862
box 18138 38862 18214 39062
use cut_M2M3_1x2 
transform 1 0 12316 0 1 38862
box 12316 38862 12392 39062
use cut_M3M4_1x2 
transform 1 0 5874 0 1 39056
box 5874 39056 5950 39256
use cut_M2M3_1x2 
transform 1 0 13396 0 1 39056
box 13396 39056 13472 39256
<< labels >>
flabel m3 s -216 35314 -140 45664 0 FreeSans 400 0 0 0 D<8>
port 6 nsew
flabel m3 s 13432 35508 13508 45690 0 FreeSans 400 0 0 0 D<3>
port 11 nsew
flabel m3 s 18472 35702 18548 45690 0 FreeSans 400 0 0 0 D<1>
port 13 nsew
flabel m3 s 10579 35896 10655 45690 0 FreeSans 400 0 0 0 D<4>
port 10 nsew
flabel m3 s 15619 36090 15695 45690 0 FreeSans 400 0 0 0 D<2>
port 12 nsew
flabel m3 s 5539 36478 5615 45690 0 FreeSans 400 0 0 0 D<6>
port 8 nsew
flabel m3 s 3352 36672 3428 45690 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8392 36866 8468 45690 0 FreeSans 400 0 0 0 D<5>
port 9 nsew
flabel m3 s 11072 50 11272 126 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew
flabel m3 s 12816 50 13016 126 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew
flabel locali s 11072 2698 11288 2758 0 FreeSans 400 0 0 0 SARN
port 3 nsew
flabel locali s 11072 1290 11288 1350 0 FreeSans 400 0 0 0 SARP
port 4 nsew
flabel locali s 20360 51744 20576 51804 0 FreeSans 400 0 0 0 DONE
port 5 nsew
flabel m3 s 20659 45690 20735 45890 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
flabel m2 s -216 40384 -16 40460 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s -232 50248 -16 50308 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 10064 498 10280 558 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel m3 s 1568 44704 1768 44904 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel m3 s 8856 0 9056 5280 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel m3 s 9648 0 9848 5280 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
<< end >>
