magic
tech sky130A
magscale 1 2
timestamp 1660667507
<< checkpaint >>
rect 0 0 1260 528
<< locali >>
rect 798 146 858 382
rect 1152 132 1368 220
rect 288 410 504 470
rect 720 146 936 206
rect 288 58 504 118
use SUNTR_PCHDL M0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_PCHDL M7
transform 1 0 0 0 1 176
box 0 176 1260 528
<< labels >>
flabel locali s 1152 132 1368 220 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 288 410 504 470 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 720 146 936 206 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 288 58 504 118 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
