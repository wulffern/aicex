magic
tech sky130A
magscale 1 2
timestamp 1658600916
<< checkpaint >>
rect 0 0 68 184
<< locali >>
rect 0 0 68 184
<< m1 >>
rect 0 0 68 184
<< viali >>
rect 6 12 62 172
<< labels >>
<< end >>
