magic
tech sky130A
magscale 1 2
timestamp 1661983200
<< checkpaint >>
rect 0 0 49444 40400
<< locali >>
rect 48676 528 48916 39872
rect 528 528 48916 768
rect 528 39632 48916 39872
rect 528 528 768 39872
rect 48676 528 48916 39872
rect 49204 0 49444 40400
rect 0 0 49444 240
rect 0 40160 49444 40400
rect 0 0 240 40400
rect 49204 0 49444 40400
rect 19432 8016 33568 8076
<< m2 >>
rect 41944 28450 42160 28510
rect 1056 1970 1272 2030
<< m1 >>
rect 30604 1056 30820 1116
use SUN_PLL_BUF xb1
transform 1 0 1056 0 1 1056
box 1056 1056 15768 12096
use SUN_PLL_LPF xb2
transform 1 0 1056 0 1 12536
box 1056 12536 41752 39344
use SUN_PLL_DIVN xc1
transform 1 0 19432 0 1 1056
box 19432 1056 33568 8092
use SUN_PLL_ROSC xd1
transform 1 0 33928 0 1 1056
box 33928 1056 40504 6464
use SUN_PLL_KICK xk1
transform 1 0 41944 0 1 1056
box 41944 1056 46000 15264
use SUN_PLL_CP xk2
transform 1 0 41944 0 1 15704
box 41944 15704 46360 26392
use SUN_PLL_PFD xk3
transform 1 0 41944 0 1 26832
box 41944 26832 46000 32592
use SUN_PLL_BIAS xl1
transform 1 0 46360 0 1 1056
box 46360 1056 48388 19776
<< labels >>
flabel locali s 48676 528 48916 39872 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 49204 0 49444 40400 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 19432 8016 33568 8076 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel m2 s 41944 28450 42160 28510 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel m1 s 30604 1056 30820 1116 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel m2 s 1056 1970 1272 2030 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
