magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 46564 39992
<< locali >>
rect 45796 528 46036 39464
rect 528 528 46036 768
rect 528 39224 46036 39464
rect 528 528 768 39464
rect 45796 528 46036 39464
rect 46324 0 46564 39992
rect 0 0 46564 240
rect 0 39752 46564 39992
rect 0 0 240 39992
rect 46324 0 46564 39992
rect 16552 8016 30688 8076
<< m2 >>
rect 39064 28450 39280 28510
rect 1056 1970 1272 2030
<< m1 >>
rect 27724 1056 27940 1116
use SUN_PLL_BUF xb1
transform 1 0 1056 0 1 1056
box 1056 1056 15768 12096
use SUN_PLL_LPF xb2
transform 1 0 1056 0 1 12536
box 1056 12536 38872 38936
use SUN_PLL_DIVN xc1
transform 1 0 16552 0 1 1056
box 16552 1056 30688 8092
use SUN_PLL_ROSC xd1
transform 1 0 31048 0 1 1056
box 31048 1056 37624 6464
use SUN_PLL_KICK xk1
transform 1 0 39064 0 1 1056
box 39064 1056 43120 15264
use SUN_PLL_CP xk2
transform 1 0 39064 0 1 15704
box 39064 15704 43480 26392
use SUN_PLL_PFD xk3
transform 1 0 39064 0 1 26832
box 39064 26832 43120 32592
use SUN_PLL_BIAS xl1
transform 1 0 43480 0 1 1056
box 43480 1056 45508 19776
<< labels >>
flabel locali s 45796 528 46036 39464 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 46324 0 46564 39992 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 16552 8016 30688 8076 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel m2 s 39064 28450 39280 28510 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel m1 s 27724 1056 27940 1116 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel m2 s 1056 1970 1272 2030 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
