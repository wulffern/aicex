** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/work/../design/SUN_PLL_SKY130NM/SUN_PLL.sch
.subckt SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U
*.ipin AVDD
*.ipin AVSS
*.ipin PWRUP_1V8
*.ipin CK_REF
*.opin CK
*.ipin IBPSR_1U
xaa0 AVDD CP_UP_N CK_REF CP_DOWN CK_FB AVSS SUN_PLL_PFD xoffset=0 yoffset=5 angle=0
xaa1 AVDD CP_UP_N VLPF CP_DOWN IBPSR_1U AVSS VLPFZ PWRUP_1V8 KICK SUN_PLL_CP xoffset=0 yoffset=5  angle=0
xaa3 AVDD KICK net1 PWRUP_1V8 AVSS PWRUP_1V8_N SUN_PLL_KICK xoffset=20 yoffset=0 angle=0
xaa4 AVDD VDD_ROSC VLPF VDD_ROSC IBPSR_1U AVSS SUN_PLL_BUF xoffset=0 yoffset=0 angle=0
xaa5 AVDD CK VDD_ROSC PWRUP_1V8 AVSS SUN_PLL_ROSC xoffset=5 yoffset=0 angle=0
xaa6 AVDD CK_FB CK PWRUP_1V8 AVSS SUN_PLL_DIVN xoffset=-310 yoffset=0 angle=0
xbb0 VLPFZ AVSS VLPF SUN_PLL_LPF xoffset=0 yoffset=5 angle=0
xbb1 IBPSR_1U PWRUP_1V8_N AVSS SUN_PLL_BIAS xoffset=5 yoffset=0 angle=0
.ends

* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_ROSC.sym # of pins=5
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_ROSC.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_ROSC.sch
.subckt SUN_PLL_ROSC  AVDD CK VDD_ROSC PWRUP_1V8 AVSS   xoffset=0 yoffset=0 angle=0
*.ipin PWRUP_1V8
*.ipin VDD_ROSC
*.ipin AVSS
*.ipin AVDD
*.opin CK
xa3 N_2 N_1 CKUP CKDWN AVDD AVSS SUN_PLL_LSCORE
xa4 CKDWN NC1 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa5 CKUP CK AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa6 AVDD AVSS SUNTR_TAPCELLB_CV xoffset=0 yoffset=0 angle=0 M=1
xb1 PWRUP_1V8 N_0 NI AVDD AVSS VDD_ROSC AVSS SUNTRB_NDX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_0 NI N_7 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_1 N_7 N_6 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_2 N_6 N_5 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_3 N_5 N_4 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_4 N_4 N_3 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_5 N_3 N_2 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_6 N_2 N_1 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb2_7 N_1 N_0 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xb3 AVDD AVSS SUNTRB_TAPCELLBAVSS_CV xoffset=0 yoffset=0 angle=0 M=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_DIVN.sym # of pins=5
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_DIVN.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_DIVN.sch
.subckt SUN_PLL_DIVN  AVDD CK_FB CK PWRUP_1V8 AVSS   xoffset=0 yoffset=0 angle=0
*.ipin PWRUP_1V8
*.ipin CK
*.ipin AVDD
*.ipin AVSS
*.opin CK_FB
xc N2 D2 PWRUP_1V8 CK_FB N2 AVDD AVSS SUNTR_DFRNQNX1_CV xoffset=0 yoffset=0 angle=0 M=1
xd N3 D3 PWRUP_1V8 D2 N3 AVDD AVSS SUNTR_DFRNQNX1_CV xoffset=0 yoffset=0 angle=0 M=1
xe N4 D4 PWRUP_1V8 D3 N4 AVDD AVSS SUNTR_DFRNQNX1_CV xoffset=0 yoffset=0 angle=0 M=1
xf N5 D5 PWRUP_1V8 D4 N5 AVDD AVSS SUNTR_DFRNQNX1_CV xoffset=0 yoffset=0 angle=0 M=1
xg N6 CK PWRUP_1V8 D5 N6 AVDD AVSS SUNTR_DFRNQNX1_CV xoffset=0 yoffset=0 angle=0 M=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_BIAS.sym # of pins=3
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BIAS.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BIAS.sch
.subckt SUN_PLL_BIAS  IBPSR_1U PWRUP_1V8_N AVSS   xoffset=0 yoffset=0 angle=0
*.ipin IBPSR_1U
*.ipin PWRUP_1V8_N
*.ipin AVSS
xa2 IBPSR_1U PWRUP_1V8_N AVSS AVSS SUNTR_NCHDL xoffset=0 yoffset=0 angle=0 M=1
xa3 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM xoffset=0 yoffset=0 angle=0 M=10
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_BUF.sym # of pins=6
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BUF.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BUF.sch
.subckt SUN_PLL_BUF  AVDD VFB VI VO VBN AVSS   xoffset=0 yoffset=0 angle=0
*.ipin AVDD
*.ipin VBN
*.ipin AVSS
*.ipin VI
*.opin VO
*.ipin VFB
xa1 VS VBN AVSS AVSS SUNTR_NCHDLCM xoffset=0 yoffset=0 angle=0 M=1
xa2 VDP VFB VS AVSS SUNTR_NCHDLA xoffset=0 yoffset=0 angle=0 M=1
xa4 VGP VI VS AVSS SUNTR_NCHDLA xoffset=0 yoffset=0 angle=0 M=1
xc1 VGP VDP AVDD AVDD SUNTR_PCHDLA xoffset=5 yoffset=0 angle=0 M=1
xc2 VDP VDP AVDD AVDD SUNTR_PCHDLA xoffset=0 yoffset=0 angle=0 M=1
xc3_0 VO VGP AVDD AVDD SUNTR_PCHDLA xoffset=0 yoffset=0 angle=0 M=1
xc3_1 VO VGP AVDD AVDD SUNTR_PCHDLA xoffset=0 yoffset=0 angle=0 M=1
xc3_2 VO VGP AVDD AVDD SUNTR_PCHDLA xoffset=0 yoffset=0 angle=0 M=1
xd2 VO AVSS SUNSAR_CAP_BSSW_CV xoffset=2 yoffset=0 angle=0 M=1
xd3 VO AVSS SUNSAR_CAP_BSSW_CV xoffset=0 yoffset=0 angle=0 M=8
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_LPF.sym # of pins=3
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LPF.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LPF.sch
.subckt SUN_PLL_LPF  VLPFZ AVSS VLPF   xoffset=0 yoffset=0 angle=0
*.ipin VLPF
*.ipin AVSS
*.ipin VLPFZ
xa1 VN5 VLPF AVSS SUNTR_RPPO8 xoffset=0 yoffset=2 angle=0 M=1
xa2 VN4 VN5 AVSS SUNTR_RPPO8 xoffset=0 yoffset=2 angle=0 M=1
xa3 VN3 VN4 AVSS SUNTR_RPPO8 xoffset=0 yoffset=2 angle=0 M=1
xa4 VN2 VN3 AVSS SUNTR_RPPO8 xoffset=0 yoffset=2 angle=0 M=1
xa5 VLPFZ VN2 AVSS SUNTR_RPPO8 xoffset=0 yoffset=2 angle=0 M=1
xb1 VLPF AVSS CAP_LPF xoffset=0 yoffset=0 angle=0 M=1
xb2 VLPF AVSS CAP_LPF xoffset=0 yoffset=0 angle=0 M=2
xb3 VLPFZ AVSS CAP_LPF xoffset=0 yoffset=0 angle=0 M=48
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_CP.sym # of pins=9
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_CP.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_CP.sch
.subckt SUN_PLL_CP  AVDD CP_UP_N LPF CP_DOWN VBN AVSS LPFZ PWRUP_1V8 KICK   xoffset=0 yoffset=0  angle=0
*.ipin AVDD
*.ipin CP_UP_N
*.ipin CP_DOWN
*.ipin VBN
*.ipin AVSS
*.opin LPF
*.ipin PWRUP_1V8
*.opin LPFZ
*.ipin KICK
xa1 VBP VBN AVSS AVSS SUNTR_NCHDLCM xoffset=0 yoffset=0 angle=0 M=1
xa2 VNS VBN AVSS AVSS SUNTR_NCHDLCM xoffset=0 yoffset=0 angle=0 M=1
xa3 LPF CP_DOWN VNS AVSS SUNTR_NCHDL xoffset=0 yoffset=0 angle=0 M=1
xa4 LPFZ KICK AVSS AVSS SUNTR_NCHDLA xoffset=0 yoffset=0 angle=0 M=10
xb1 VBP VBP AVDD AVDD SUNTR_PCHDLCM xoffset=5 yoffset=0 angle=0 M=1
xb2 VPS VBP AVDD AVDD SUNTR_PCHDLCM xoffset=0 yoffset=0 angle=0 M=1
xb3 LPF CP_UP_N VPS AVDD SUNTR_PCHDL xoffset=0 yoffset=0 angle=0 M=1
xb4 LPF PWRUP_1V8 AVDD AVDD SUNTR_PCHDL xoffset=0 yoffset=0 angle=0 M=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_PFD.sym # of pins=6
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_PFD.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_PFD.sch
.subckt SUN_PLL_PFD  AVDD CP_UP_N CK_REF CP_DOWN CK_FB AVSS   xoffset=0 yoffset=0 angle=0
*.ipin CK_FB
*.ipin CK_REF
*.opin CP_UP_N
*.opin CP_DOWN
*.ipin AVDD
*.ipin AVSS
xa0 AVDD AVSS SUNTR_TAPCELLB_CV xoffset=0 yoffset=0 angle=0 M=1
xa1 CFB CK_REF CP_DUP_N AVDD AVSS SUNTR_DFTSPCX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa2 CP_DUP_N CP_UP AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa2a CP_UP CP_UP_N AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa3 CP_DUP_N CP_DOWN_N CFB AVDD AVSS SUNTR_NRX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa5 CFB CK_FB CP_DOWN_N AVDD AVSS SUNTR_DFTSPCX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa6 CP_DOWN_N CP_DOWN AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_KICK.sym # of pins=6
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_KICK.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_KICK.sch
.subckt SUN_PLL_KICK  AVDD KICK KICK_N PWRUP_1V8 AVSS PWRUP_1V8_N   xoffset=0 yoffset=0 angle=0
*.ipin PWRUP_1V8
*.opin KICK
*.opin KICK_N
*.ipin AVDD
*.ipin AVSS
*.opin PWRUP_1V8_N
xa1a AVDD AVSS SUNTR_TAPCELLB_CV xoffset=0 yoffset=0 angle=0 M=1
xa1b PWRUP_1V8 PWRUP_1V8_N AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa1c PWRUP_1V8_N N1 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa1capd AVSS N1 SUNTR_DCAPX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa2 N1 N2 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa3a N2 N3 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa3capb AVSS N3 SUNTR_DCAPX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa4 N3 N4 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa5a N4 N5 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa5capb AVSS N5 SUNTR_DCAPX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa6 N5 N6 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa7 N6 N7 AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa8 PWRUP_1V8_N N7 KICK AVDD AVSS SUNTR_NRX1_CV xoffset=0 yoffset=0 angle=0 M=1
xa9 KICK KICK_N AVDD AVSS SUNTR_IVX1_CV xoffset=0 yoffset=0 angle=0 M=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sym # of pins=6
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sch
.subckt SUN_PLL_LSCORE  A AN YN Y AVDD AVSS
*.ipin AVDD
*.ipin A
*.ipin AN
*.opin Y
*.opin YN
*.ipin AVSS
xb1_0 Y AN AVSS AVSS SUNTR_NCHDL xoffset=0 yoffset=0 angle=0 M=1
xb1_1 Y AN AVSS AVSS SUNTR_NCHDL xoffset=0 yoffset=0 angle=0 M=1
xb2_0 YN A AVSS AVSS SUNTR_NCHDL xoffset=0 yoffset=0 angle=0 M=1
xb2_1 YN A AVSS AVSS SUNTR_NCHDL xoffset=0 yoffset=0 angle=0 M=1
xc1a net2 YN AVDD AVDD SUNTR_PCHDL xoffset=0 yoffset=0 angle=0 M=1
xc1b Y YN net2 AVDD SUNTR_PCHDL xoffset=0 yoffset=0 angle=0 M=1
xc2a net1 Y AVDD AVDD SUNTR_PCHDL xoffset=0 yoffset=0 angle=0 M=1
xc2b YN Y net1 AVDD SUNTR_PCHDL xoffset=0 yoffset=0 angle=0 M=1
.ends


* expanding   symbol:  SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV.sym # of pins=2
** sym_path:
*+ /Users/wulff/prog/aicex/ip/sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV.sym
** sch_path:
*+ /Users/wulff/prog/aicex/ip/sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV.sch
.subckt SUNSAR_CAP_BSSW_CV  A B   xoffset=0 yoffset=0 angle=0 M=1
*.iopin A
*.iopin B
R1 A NC0 sky130_fd_pr__res_generic_m1 W=0.44 L=0.36 m=1
R2 B NC1 sky130_fd_pr__res_generic_m1 W=0.44 L=0.36 m=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/CAP_LPF.sym # of pins=2
** sym_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/CAP_LPF.sym
** sch_path: /Users/wulff/prog/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/CAP_LPF.sch
.subckt CAP_LPF  A B   xoffset=0 yoffset=0 angle=0 M=1
*.iopin A
*.iopin B
R1 A NC0 sky130_fd_pr__res_generic_m3 W=0.4 L=0.4 m=1
R2 B NC1 sky130_fd_pr__res_generic_m3 W=0.4 L=0.4 m=1
.ends

.end
