magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 960
<< locali >>
rect 800 850 968 910
rect 968 850 1520 910
rect 968 850 1028 910
rect 1890 130 1950 830
rect 770 210 830 430
rect 770 530 830 750
rect 1490 210 1550 430
rect 1490 530 1550 750
<< m3 >>
rect 1400 0 1600 960
rect 680 0 880 960
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1160 960
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL MP2
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use cut_M1M4_2x1 
transform 1 0 1400 0 1 50
box 1400 50 1600 118
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
<< labels >>
flabel locali s 2200 120 2440 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -120 120 120 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel locali s 1800 770 2040 830 0 FreeSans 400 0 0 0 RST_N
port 4 nsew
flabel locali s 280 770 520 830 0 FreeSans 400 0 0 0 EN
port 5 nsew
flabel locali s 280 450 520 510 0 FreeSans 400 0 0 0 LCK_N
port 6 nsew
flabel locali s 680 850 920 910 0 FreeSans 400 0 0 0 CHL
port 7 nsew
flabel m3 s 1400 0 1600 960 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 680 0 880 960 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
