magic
tech sky130A
magscale 1 2
timestamp 1660916687
<< checkpaint >>
rect -1560 -1920 46660 54640
<< locali >>
rect 45892 -1392 46132 54112
rect -1032 -1392 46132 -1152
rect -1032 53872 46132 54112
rect -1032 -1392 -792 54112
rect 45892 -1392 46132 54112
rect 46420 -1920 46660 54640
rect -1560 -1920 46660 -1680
rect -1560 54400 46660 54640
rect -1560 -1920 -1320 54640
rect 46420 -1920 46660 54640
rect 15376 7248 29512 7308
rect 38620 26626 38836 26686
rect 26548 1554 26764 1614
rect 684 146 900 206
use SUN_PLL_BUF xb1
transform 1 0 360 0 1 0
box 360 0 15072 23712
use SUN_PLL_LPF xb2
transform 1 0 360 0 1 24592
box 360 24592 39904 52720
use SUN_PLL_DIVN xc1
transform 1 0 16144 0 1 1056
box 16144 1056 30280 8076
use SUN_PLL_ROSC xd1
transform 1 0 30280 0 1 0
box 30280 0 36856 5408
use SUN_PLL_KICK xk1
transform 1 0 38296 0 1 0
box 38296 0 42352 14208
use SUN_PLL_CP xk2
transform 1 0 38296 0 1 15088
box 38296 15088 42712 25776
use SUN_PLL_PFD xk3
transform 1 0 38296 0 1 25776
box 38296 25776 42352 31536
use SUN_PLL_BIAS xl1
transform 1 0 42712 0 1 0
box 42712 0 44740 18720
<< labels >>
flabel locali s 45892 -1392 46132 54112 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 46420 -1920 46660 54640 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 15376 7248 29512 7308 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel locali s 38620 26626 38836 26686 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel locali s 26548 1554 26764 1614 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel locali s 684 146 900 206 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
