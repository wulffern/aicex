magic
tech sky130A
magscale 1 2
timestamp 1658699483
<< checkpaint >>
rect 0 0 76 200
<< m3 >>
rect 0 0 76 200
<< m4 >>
rect 0 0 76 200
<< v3 >>
rect 6 12 70 188
<< labels >>
<< end >>
