magic
tech sky130A
magscale 1 2
timestamp 1660667507
<< checkpaint >>
rect -640 -640 1720 3500
<< locali >>
rect -640 -640 1720 -528
rect -640 -640 1720 -528
rect -640 -640 -528 3500
rect -640 3388 1720 3500
rect 1608 -640 1720 3500
rect -640 -640 1720 -528
rect 810 2750 1134 2970
rect -54 2750 270 2970
<< ptapc >>
rect -620 -640 -540 -560
rect -540 -640 -460 -560
rect -460 -640 -380 -560
rect -380 -640 -300 -560
rect -300 -640 -220 -560
rect -220 -640 -140 -560
rect -140 -640 -60 -560
rect -60 -640 20 -560
rect 20 -640 100 -560
rect 100 -640 180 -560
rect 180 -640 260 -560
rect 260 -640 340 -560
rect 340 -640 420 -560
rect 420 -640 500 -560
rect 500 -640 580 -560
rect 580 -640 660 -560
rect 660 -640 740 -560
rect 740 -640 820 -560
rect 820 -640 900 -560
rect 900 -640 980 -560
rect 980 -640 1060 -560
rect 1060 -640 1140 -560
rect 1140 -640 1220 -560
rect 1220 -640 1300 -560
rect 1300 -640 1380 -560
rect 1380 -640 1460 -560
rect 1460 -640 1540 -560
rect 1540 -640 1620 -560
rect 1620 -640 1700 -560
rect -640 -610 -560 -530
rect -640 -530 -560 -450
rect -640 -450 -560 -370
rect -640 -370 -560 -290
rect -640 -290 -560 -210
rect -640 -210 -560 -130
rect -640 -130 -560 -50
rect -640 -50 -560 30
rect -640 30 -560 110
rect -640 110 -560 190
rect -640 190 -560 270
rect -640 270 -560 350
rect -640 350 -560 430
rect -640 430 -560 510
rect -640 510 -560 590
rect -640 590 -560 670
rect -640 670 -560 750
rect -640 750 -560 830
rect -640 830 -560 910
rect -640 910 -560 990
rect -640 990 -560 1070
rect -640 1070 -560 1150
rect -640 1150 -560 1230
rect -640 1230 -560 1310
rect -640 1310 -560 1390
rect -640 1390 -560 1470
rect -640 1470 -560 1550
rect -640 1550 -560 1630
rect -640 1630 -560 1710
rect -640 1710 -560 1790
rect -640 1790 -560 1870
rect -640 1870 -560 1950
rect -640 1950 -560 2030
rect -640 2030 -560 2110
rect -640 2110 -560 2190
rect -640 2190 -560 2270
rect -640 2270 -560 2350
rect -640 2350 -560 2430
rect -640 2430 -560 2510
rect -640 2510 -560 2590
rect -640 2590 -560 2670
rect -640 2670 -560 2750
rect -640 2750 -560 2830
rect -640 2830 -560 2910
rect -640 2910 -560 2990
rect -640 2990 -560 3070
rect -640 3070 -560 3150
rect -640 3150 -560 3230
rect -640 3230 -560 3310
rect -640 3310 -560 3390
rect -640 3390 -560 3470
rect -620 3388 -540 3468
rect -540 3388 -460 3468
rect -460 3388 -380 3468
rect -380 3388 -300 3468
rect -300 3388 -220 3468
rect -220 3388 -140 3468
rect -140 3388 -60 3468
rect -60 3388 20 3468
rect 20 3388 100 3468
rect 100 3388 180 3468
rect 180 3388 260 3468
rect 260 3388 340 3468
rect 340 3388 420 3468
rect 420 3388 500 3468
rect 500 3388 580 3468
rect 580 3388 660 3468
rect 660 3388 740 3468
rect 740 3388 820 3468
rect 820 3388 900 3468
rect 900 3388 980 3468
rect 980 3388 1060 3468
rect 1060 3388 1140 3468
rect 1140 3388 1220 3468
rect 1220 3388 1300 3468
rect 1300 3388 1380 3468
rect 1380 3388 1460 3468
rect 1460 3388 1540 3468
rect 1540 3388 1620 3468
rect 1620 3388 1700 3468
rect 1608 -610 1688 -530
rect 1608 -530 1688 -450
rect 1608 -450 1688 -370
rect 1608 -370 1688 -290
rect 1608 -290 1688 -210
rect 1608 -210 1688 -130
rect 1608 -130 1688 -50
rect 1608 -50 1688 30
rect 1608 30 1688 110
rect 1608 110 1688 190
rect 1608 190 1688 270
rect 1608 270 1688 350
rect 1608 350 1688 430
rect 1608 430 1688 510
rect 1608 510 1688 590
rect 1608 590 1688 670
rect 1608 670 1688 750
rect 1608 750 1688 830
rect 1608 830 1688 910
rect 1608 910 1688 990
rect 1608 990 1688 1070
rect 1608 1070 1688 1150
rect 1608 1150 1688 1230
rect 1608 1230 1688 1310
rect 1608 1310 1688 1390
rect 1608 1390 1688 1470
rect 1608 1470 1688 1550
rect 1608 1550 1688 1630
rect 1608 1630 1688 1710
rect 1608 1710 1688 1790
rect 1608 1790 1688 1870
rect 1608 1870 1688 1950
rect 1608 1950 1688 2030
rect 1608 2030 1688 2110
rect 1608 2110 1688 2190
rect 1608 2190 1688 2270
rect 1608 2270 1688 2350
rect 1608 2350 1688 2430
rect 1608 2430 1688 2510
rect 1608 2510 1688 2590
rect 1608 2590 1688 2670
rect 1608 2670 1688 2750
rect 1608 2750 1688 2830
rect 1608 2830 1688 2910
rect 1608 2910 1688 2990
rect 1608 2990 1688 3070
rect 1608 3070 1688 3150
rect 1608 3150 1688 3230
rect 1608 3230 1688 3310
rect 1608 3310 1688 3390
rect 1608 3390 1688 3470
<< ptap >>
rect -640 -640 1720 -528
rect -640 -640 -528 3500
rect -640 3388 1720 3500
rect 1608 -640 1720 3500
use SUNTR_RES25 XA1
transform 1 0 0 0 1 0
box 0 0 1080 2860
<< labels >>
flabel locali s -640 -640 1720 -528 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 810 2750 1134 2970 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s -54 2750 270 2970 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
