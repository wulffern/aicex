magic
tech sky130A
magscale 1 2
timestamp 1658775803
<< checkpaint >>
rect 0 0 2520 11616
<< locali >>
rect 432 5074 600 5134
rect 600 4458 864 4518
rect 600 4458 660 5134
rect 432 6482 600 6542
rect 600 5866 864 5926
rect 600 5866 660 6542
rect 1860 4370 2088 4430
rect 1656 4106 1860 4166
rect 1860 4106 1920 4430
rect 432 8946 600 9006
rect 600 8682 864 8742
rect 600 8682 660 9006
rect 402 8946 462 9358
rect 480 9942 600 10002
rect 600 9738 864 9798
rect 600 9738 660 10002
rect 480 10002 540 10062
rect 480 10294 600 10354
rect 600 10090 864 10150
rect 600 10090 660 10354
rect 480 10354 540 10414
rect 432 11058 600 11118
rect 600 10618 864 10678
rect 600 10618 660 11118
rect 1656 6570 1824 6630
rect 1824 7186 2088 7246
rect 1824 6570 1884 7246
rect 1980 4018 2196 4078
rect 324 3314 540 3374
rect 324 10706 540 10766
rect 1548 11146 1764 11206
rect 324 7538 540 7598
rect 756 9034 972 9094
<< m1 >>
rect 432 5778 600 5838
rect 600 3050 864 3110
rect 600 3050 660 5846
rect 2088 8594 2256 8654
rect 1656 762 2256 822
rect 2256 762 2316 8662
rect 432 9650 600 9710
rect 600 8330 864 8390
rect 600 8330 660 9718
rect 1656 5162 1824 5222
rect 1824 7890 2088 7950
rect 1824 5162 1884 7958
<< m3 >>
rect 2186 4810 2262 7122
rect 340 5066 540 5142
rect 1055 5092 1131 5292
rect 1215 5796 1291 5996
rect 1390 6500 1466 6700
rect 2124 4810 2324 5010
rect 1548 0 1748 11616
rect 756 0 956 11616
rect 1548 0 1748 11616
rect 756 0 956 11616
<< m2 >>
rect 340 2250 540 2326
rect 340 490 540 566
rect 1564 754 1764 830
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use SARMRYX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2520 4224
use SWX2_CV XA2
transform 1 0 0 0 1 4224
box 0 4224 2520 4928
use SWX2_CV XA3
transform 1 0 0 0 1 4928
box 0 4928 2520 5632
use SWX2_CV XA4
transform 1 0 0 0 1 5632
box 0 5632 2520 6336
use SWX2_CV XA5
transform 1 0 0 0 1 6336
box 0 6336 2520 7040
use SARCEX1_CV XA6
transform 1 0 0 0 1 7040
box 0 7040 2520 8448
use IVX1_CV XA7
transform 1 0 0 0 1 8448
box 0 8448 2520 8800
use IVX1_CV XA8
transform 1 0 0 0 1 8800
box 0 8800 2520 9152
use NDX1_CV XA9
transform 1 0 0 0 1 9152
box 0 9152 2520 9856
use IVX1_CV XA10
transform 1 0 0 0 1 9856
box 0 9856 2520 10208
use NRX1_CV XA11
transform 1 0 0 0 1 10208
box 0 10208 2520 10912
use IVX1_CV XA12
transform 1 0 0 0 1 10912
box 0 10912 2520 11264
use TAPCELLB_CV XA13
transform 1 0 0 0 1 11264
box 0 11264 2520 11616
use DMY_CV XA14
transform 1 0 0 0 1 11616
box 0 11616 0 11616
use cut_M1M2_2x1 
transform 1 0 324 0 1 5778
box 324 5778 508 5846
use cut_M1M2_2x1 
transform 1 0 756 0 1 3050
box 756 3050 940 3118
use cut_M1M2_2x1 
transform 1 0 1980 0 1 8594
box 1980 8594 2164 8662
use cut_M1M2_2x1 
transform 1 0 1548 0 1 762
box 1548 762 1732 830
use cut_M1M2_2x1 
transform 1 0 324 0 1 9650
box 324 9650 508 9718
use cut_M1M2_2x1 
transform 1 0 756 0 1 8330
box 756 8330 940 8398
use cut_M1M2_2x1 
transform 1 0 1548 0 1 5162
box 1548 5162 1732 5230
use cut_M1M2_2x1 
transform 1 0 1980 0 1 7890
box 1980 7890 2164 7958
use cut_M1M4_2x1 
transform 1 0 340 0 1 5066
box 340 5066 540 5142
use cut_M1M4_1x2 
transform 1 0 1055 0 1 5092
box 1055 5092 1131 5292
use cut_M1M4_1x2 
transform 1 0 1215 0 1 5796
box 1215 5796 1291 5996
use cut_M1M4_1x2 
transform 1 0 1390 0 1 6500
box 1390 6500 1466 6700
use cut_M2M3_2x1 
transform 1 0 1564 0 1 754
box 1564 754 1764 830
use cut_M2M3_2x1 
transform 1 0 340 0 1 490
box 340 490 540 566
use cut_M2M3_2x1 
transform 1 0 340 0 1 490
box 340 490 540 566
use cut_M2M3_2x1 
transform 1 0 340 0 1 2250
box 340 2250 540 2326
use cut_M2M3_2x1 
transform 1 0 340 0 1 2250
box 340 2250 540 2326
<< labels >>
flabel m2 s 340 2250 540 2326 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1980 4018 2196 4078 0 FreeSans 400 0 0 0 RST_N
port 4 nsew
flabel m2 s 340 490 540 566 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 324 3314 540 3374 0 FreeSans 400 0 0 0 CMP_ON
port 2 nsew
flabel m2 s 1564 754 1764 830 0 FreeSans 400 0 0 0 ENO
port 5 nsew
flabel m3 s 340 5066 540 5142 0 FreeSans 400 0 0 0 CN1
port 10 nsew
flabel m3 s 1055 5092 1131 5292 0 FreeSans 400 0 0 0 CP1
port 8 nsew
flabel m3 s 1215 5796 1291 5996 0 FreeSans 400 0 0 0 CP0
port 7 nsew
flabel m3 s 1390 6500 1466 6700 0 FreeSans 400 0 0 0 CN0
port 9 nsew
flabel locali s 324 10706 540 10766 0 FreeSans 400 0 0 0 CEIN
port 11 nsew
flabel locali s 1548 11146 1764 11206 0 FreeSans 400 0 0 0 CEO
port 12 nsew
flabel locali s 324 7538 540 7598 0 FreeSans 400 0 0 0 CKS
port 13 nsew
flabel locali s 756 9034 972 9094 0 FreeSans 400 0 0 0 DONE
port 6 nsew
flabel m3 s 2124 4810 2324 5010 0 FreeSans 400 0 0 0 VREF
port 14 nsew
flabel m3 s 1548 0 1748 11616 0 FreeSans 400 0 0 0 AVDD
port 15 nsew
flabel m3 s 756 0 956 11616 0 FreeSans 400 0 0 0 AVSS
port 16 nsew
<< end >>
