magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 640
<< locali >>
rect 720 210 874 270
rect 720 370 874 430
rect 874 210 1380 270
rect 874 370 1380 430
rect 874 210 934 430
rect 330 130 390 510
rect 1710 130 1770 510
rect 270 130 450 190
rect 630 210 810 270
rect 2010 120 2190 200
rect -90 120 90 200
<< poly >>
rect 270 142 1830 178
rect 270 462 1830 498
<< m2 >>
rect 1380 50 1534 118
rect 1380 530 1534 598
rect 1534 530 1862 598
rect 1534 50 1602 598
<< m3 >>
rect 1770 530 1954 714
rect 630 0 814 640
rect 630 0 814 640
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use cut_M3M4_2x2 
transform 1 0 1770 0 1 530
box 1770 530 1954 714
use cut_M1M3_2x1 
transform 1 0 1290 0 1 50
box 1290 50 1474 118
use cut_M1M3_2x1 
transform 1 0 1290 0 1 530
box 1290 530 1474 598
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
<< labels >>
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 630 210 810 270 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 3 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 4 nsew
flabel m3 s 1770 530 1954 714 0 FreeSans 400 0 0 0 VREF
port 5 nsew
flabel m3 s 630 0 814 640 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
