magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 1280
<< locali >>
rect 1350 530 1410 750
rect 1350 850 1410 1070
rect 720 210 874 270
rect 720 530 874 590
rect 720 690 874 750
rect 874 210 934 750
rect 1166 370 1380 430
rect 720 1170 1166 1230
rect 1166 370 1226 1230
rect 1380 50 1534 110
rect 1534 1090 1740 1150
rect 1534 50 1594 1150
rect 630 50 1470 110
rect 2010 120 2190 200
rect -90 120 90 200
rect 270 770 450 830
rect 270 450 450 510
rect 1650 130 1830 190
rect 270 130 450 190
rect 1290 370 1470 430
<< poly >>
rect 270 462 1830 498
rect 270 782 1830 818
rect 270 1102 1830 1138
<< m3 >>
rect 1290 0 1474 1280
rect 630 0 814 1280
rect 1290 0 1474 1280
rect 630 0 814 1280
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1050 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1050 1280
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL MP2
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use PCHDL MP3
transform 1 0 1050 0 1 960
box 1050 960 2100 1280
use cut_M1M4_2x1 
transform 1 0 1290 0 1 210
box 1290 210 1474 278
use cut_M1M4_2x1 
transform 1 0 1290 0 1 1170
box 1290 1170 1474 1238
use cut_M1M4_2x1 
transform 1 0 630 0 1 370
box 630 370 814 438
use cut_M1M4_2x1 
transform 1 0 630 0 1 850
box 630 850 814 918
use cut_M1M4_2x1 
transform 1 0 630 0 1 1010
box 630 1010 814 1078
<< labels >>
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 270 770 450 830 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 1650 130 1830 190 0 FreeSans 400 0 0 0 RST_N
port 5 nsew
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 EN
port 6 nsew
flabel locali s 1290 370 1470 430 0 FreeSans 400 0 0 0 ENO
port 7 nsew
flabel m3 s 1290 0 1474 1280 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 1280 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
