magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 39832 49848
<< locali >>
rect 39532 0 39832 49848
rect 0 0 39832 300
rect 0 49548 39832 49848
rect 0 0 300 49848
rect 39532 0 39832 49848
rect 300 636 460 748
rect 300 5048 460 5160
rect 300 9460 460 9572
rect 300 13872 460 13984
rect 300 18284 460 18396
rect 4516 21706 5092 21926
rect 1060 4058 1636 4278
<< m3 >>
rect 22400 0 22616 484
rect 39268 404 39608 480
rect 39268 1364 39608 1440
rect 39268 2324 39608 2400
rect 39268 3284 39608 3360
rect 39268 4244 39608 4320
rect 39268 5204 39608 5280
rect 39268 6164 39608 6240
rect 39268 7124 39608 7200
rect 39268 8084 39608 8160
rect 39268 9044 39608 9120
rect 39268 10004 39608 10080
rect 39268 10964 39608 11040
rect 39268 11924 39608 12000
rect 39268 12884 39608 12960
rect 39268 13844 39608 13920
rect 39268 14804 39608 14880
rect 39268 15764 39608 15840
rect 39268 16724 39608 16800
rect 39268 17684 39608 17760
rect 39268 18644 39608 18720
rect 39268 19604 39608 19680
rect 39268 20564 39608 20640
rect 39268 21524 39608 21600
rect 39268 22484 39608 22560
rect 39268 23444 39608 23520
rect 39268 24404 39608 24480
rect 39268 25364 39608 25440
rect 39268 26324 39608 26400
rect 39268 27284 39608 27360
rect 39268 28244 39608 28320
rect 39268 29204 39608 29280
rect 39268 30164 39608 30240
rect 39268 31124 39608 31200
rect 39268 32084 39608 32160
rect 39268 33044 39608 33120
rect 39268 34004 39608 34080
rect 39268 34964 39608 35040
rect 39268 35924 39608 36000
rect 39268 36884 39608 36960
rect 39268 37844 39608 37920
rect 39268 38804 39608 38880
rect 39268 39764 39608 39840
rect 39268 40724 39608 40800
rect 39268 41684 39608 41760
rect 39268 42644 39608 42720
rect 39268 43604 39608 43680
rect 39268 44564 39608 44640
rect 39268 45524 39608 45600
rect 39268 46484 39608 46560
rect 39268 47444 39608 47520
rect 39268 48404 39608 48480
<< m1 >>
rect 1152 8470 1364 8530
rect 1364 4058 4608 4118
rect 1364 4058 1424 8530
rect 1152 17294 1508 17354
rect 1508 12882 4608 12942
rect 1508 12882 1568 17354
rect 4608 21706 4760 21766
rect 4760 4084 5848 4144
rect 4760 5044 5848 5104
rect 4760 6004 5848 6064
rect 4760 6964 5848 7024
rect 4760 7924 5848 7984
rect 4760 8884 5848 8944
rect 4760 9844 5848 9904
rect 4760 10804 5848 10864
rect 4760 11764 5848 11824
rect 4760 12724 5848 12784
rect 4760 13684 5848 13744
rect 4760 14644 5848 14704
rect 4760 15604 5848 15664
rect 4760 16564 5848 16624
rect 4760 17524 5848 17584
rect 4760 18484 5848 18544
rect 4760 19444 5848 19504
rect 4760 20404 5848 20464
rect 4760 21364 5848 21424
rect 4760 22324 5848 22384
rect 4760 23284 5848 23344
rect 4760 24244 5848 24304
rect 4760 25204 5848 25264
rect 4760 26164 5848 26224
rect 4760 27124 5848 27184
rect 4760 28084 5848 28144
rect 4760 29044 5848 29104
rect 4760 30004 5848 30064
rect 4760 30964 5848 31024
rect 4760 31924 5848 31984
rect 4760 32884 5848 32944
rect 4760 33844 5848 33904
rect 4760 34804 5848 34864
rect 4760 35764 5848 35824
rect 4760 36724 5848 36784
rect 4760 37684 5848 37744
rect 4760 38644 5848 38704
rect 4760 39604 5848 39664
rect 4760 40564 5848 40624
rect 4760 41524 5848 41584
rect 4760 42484 5848 42544
rect 4760 43444 5848 43504
rect 4760 44404 5848 44464
rect 4760 45364 5848 45424
rect 4760 46324 5848 46384
rect 4760 47284 5848 47344
rect 4760 48244 5848 48304
rect 4760 49204 5848 49264
rect 4760 4084 4820 49264
<< m2 >>
rect 1160 12882 1388 12958
rect 1388 8470 4616 8546
rect 1388 8470 1464 12958
rect 1160 21706 1676 21782
rect 1676 17294 4616 17370
rect 1676 17294 1752 21782
rect 1160 4058 1324 4134
rect 1324 1204 5848 1280
rect 1324 2164 5848 2240
rect 1324 3124 5848 3200
rect 1324 1204 1400 4134
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa10
transform 1 0 444 0 1 620
box 444 620 5708 4856
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa20
transform 1 0 444 0 1 5032
box 444 5032 5708 9268
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa30
transform 1 0 444 0 1 9444
box 444 9444 5708 13680
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa40
transform 1 0 444 0 1 13856
box 444 13856 5708 18092
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa50
transform 1 0 444 0 1 18268
box 444 18268 5708 22504
use CAP_LPF xb10
transform -1 0 39388 0 1 444
box 39388 444 73068 1404
use CAP_LPF xb20
transform -1 0 39388 0 1 1404
box 39388 1404 73068 2364
use CAP_LPF xb21
transform -1 0 39388 0 1 2364
box 39388 2364 73068 3324
use CAP_LPF xb30
transform -1 0 39388 0 1 3324
box 39388 3324 73068 4284
use CAP_LPF xb31
transform -1 0 39388 0 1 4284
box 39388 4284 73068 5244
use CAP_LPF xb32
transform -1 0 39388 0 1 5244
box 39388 5244 73068 6204
use CAP_LPF xb33
transform -1 0 39388 0 1 6204
box 39388 6204 73068 7164
use CAP_LPF xb34
transform -1 0 39388 0 1 7164
box 39388 7164 73068 8124
use CAP_LPF xb35
transform -1 0 39388 0 1 8124
box 39388 8124 73068 9084
use CAP_LPF xb36
transform -1 0 39388 0 1 9084
box 39388 9084 73068 10044
use CAP_LPF xb37
transform -1 0 39388 0 1 10044
box 39388 10044 73068 11004
use CAP_LPF xb38
transform -1 0 39388 0 1 11004
box 39388 11004 73068 11964
use CAP_LPF xb39
transform -1 0 39388 0 1 11964
box 39388 11964 73068 12924
use CAP_LPF xb310
transform -1 0 39388 0 1 12924
box 39388 12924 73068 13884
use CAP_LPF xb311
transform -1 0 39388 0 1 13884
box 39388 13884 73068 14844
use CAP_LPF xb312
transform -1 0 39388 0 1 14844
box 39388 14844 73068 15804
use CAP_LPF xb313
transform -1 0 39388 0 1 15804
box 39388 15804 73068 16764
use CAP_LPF xb314
transform -1 0 39388 0 1 16764
box 39388 16764 73068 17724
use CAP_LPF xb315
transform -1 0 39388 0 1 17724
box 39388 17724 73068 18684
use CAP_LPF xb316
transform -1 0 39388 0 1 18684
box 39388 18684 73068 19644
use CAP_LPF xb317
transform -1 0 39388 0 1 19644
box 39388 19644 73068 20604
use CAP_LPF xb318
transform -1 0 39388 0 1 20604
box 39388 20604 73068 21564
use CAP_LPF xb319
transform -1 0 39388 0 1 21564
box 39388 21564 73068 22524
use CAP_LPF xb320
transform -1 0 39388 0 1 22524
box 39388 22524 73068 23484
use CAP_LPF xb321
transform -1 0 39388 0 1 23484
box 39388 23484 73068 24444
use CAP_LPF xb322
transform -1 0 39388 0 1 24444
box 39388 24444 73068 25404
use CAP_LPF xb323
transform -1 0 39388 0 1 25404
box 39388 25404 73068 26364
use CAP_LPF xb324
transform -1 0 39388 0 1 26364
box 39388 26364 73068 27324
use CAP_LPF xb325
transform -1 0 39388 0 1 27324
box 39388 27324 73068 28284
use CAP_LPF xb326
transform -1 0 39388 0 1 28284
box 39388 28284 73068 29244
use CAP_LPF xb327
transform -1 0 39388 0 1 29244
box 39388 29244 73068 30204
use CAP_LPF xb328
transform -1 0 39388 0 1 30204
box 39388 30204 73068 31164
use CAP_LPF xb329
transform -1 0 39388 0 1 31164
box 39388 31164 73068 32124
use CAP_LPF xb330
transform -1 0 39388 0 1 32124
box 39388 32124 73068 33084
use CAP_LPF xb331
transform -1 0 39388 0 1 33084
box 39388 33084 73068 34044
use CAP_LPF xb332
transform -1 0 39388 0 1 34044
box 39388 34044 73068 35004
use CAP_LPF xb333
transform -1 0 39388 0 1 35004
box 39388 35004 73068 35964
use CAP_LPF xb334
transform -1 0 39388 0 1 35964
box 39388 35964 73068 36924
use CAP_LPF xb335
transform -1 0 39388 0 1 36924
box 39388 36924 73068 37884
use CAP_LPF xb336
transform -1 0 39388 0 1 37884
box 39388 37884 73068 38844
use CAP_LPF xb337
transform -1 0 39388 0 1 38844
box 39388 38844 73068 39804
use CAP_LPF xb338
transform -1 0 39388 0 1 39804
box 39388 39804 73068 40764
use CAP_LPF xb339
transform -1 0 39388 0 1 40764
box 39388 40764 73068 41724
use CAP_LPF xb340
transform -1 0 39388 0 1 41724
box 39388 41724 73068 42684
use CAP_LPF xb341
transform -1 0 39388 0 1 42684
box 39388 42684 73068 43644
use CAP_LPF xb342
transform -1 0 39388 0 1 43644
box 39388 43644 73068 44604
use CAP_LPF xb343
transform -1 0 39388 0 1 44604
box 39388 44604 73068 45564
use CAP_LPF xb344
transform -1 0 39388 0 1 45564
box 39388 45564 73068 46524
use CAP_LPF xb345
transform -1 0 39388 0 1 46524
box 39388 46524 73068 47484
use CAP_LPF xb346
transform -1 0 39388 0 1 47484
box 39388 47484 73068 48444
use CAP_LPF xb347
transform -1 0 39388 0 1 48444
box 39388 48444 73068 49404
use cut_M1M4_2x1 
transform 1 0 22408 0 1 0
box 22408 0 22608 76
use cut_M1M2_2x1 
transform 1 0 1060 0 1 8470
box 1060 8470 1244 8538
use cut_M1M2_2x1 
transform 1 0 4516 0 1 4058
box 4516 4058 4700 4126
use cut_M1M3_2x1 
transform 1 0 1060 0 1 12882
box 1060 12882 1260 12958
use cut_M1M3_2x1 
transform 1 0 4516 0 1 8470
box 4516 8470 4716 8546
use cut_M1M2_2x1 
transform 1 0 1060 0 1 17294
box 1060 17294 1244 17362
use cut_M1M2_2x1 
transform 1 0 4516 0 1 12882
box 4516 12882 4700 12950
use cut_M1M3_2x1 
transform 1 0 1060 0 1 21706
box 1060 21706 1260 21782
use cut_M1M3_2x1 
transform 1 0 4516 0 1 17294
box 4516 17294 4716 17370
use cut_M1M2_2x1 
transform 1 0 4516 0 1 21706
box 4516 21706 4700 21774
use cut_M2M4_2x1 
transform 1 0 5748 0 1 4084
box 5748 4084 5948 4160
use cut_M2M4_2x1 
transform 1 0 5748 0 1 5044
box 5748 5044 5948 5120
use cut_M2M4_2x1 
transform 1 0 5748 0 1 6004
box 5748 6004 5948 6080
use cut_M2M4_2x1 
transform 1 0 5748 0 1 6964
box 5748 6964 5948 7040
use cut_M2M4_2x1 
transform 1 0 5748 0 1 7924
box 5748 7924 5948 8000
use cut_M2M4_2x1 
transform 1 0 5748 0 1 8884
box 5748 8884 5948 8960
use cut_M2M4_2x1 
transform 1 0 5748 0 1 9844
box 5748 9844 5948 9920
use cut_M2M4_2x1 
transform 1 0 5748 0 1 10804
box 5748 10804 5948 10880
use cut_M2M4_2x1 
transform 1 0 5748 0 1 11764
box 5748 11764 5948 11840
use cut_M2M4_2x1 
transform 1 0 5748 0 1 12724
box 5748 12724 5948 12800
use cut_M2M4_2x1 
transform 1 0 5748 0 1 13684
box 5748 13684 5948 13760
use cut_M2M4_2x1 
transform 1 0 5748 0 1 14644
box 5748 14644 5948 14720
use cut_M2M4_2x1 
transform 1 0 5748 0 1 15604
box 5748 15604 5948 15680
use cut_M2M4_2x1 
transform 1 0 5748 0 1 16564
box 5748 16564 5948 16640
use cut_M2M4_2x1 
transform 1 0 5748 0 1 17524
box 5748 17524 5948 17600
use cut_M2M4_2x1 
transform 1 0 5748 0 1 18484
box 5748 18484 5948 18560
use cut_M2M4_2x1 
transform 1 0 5748 0 1 19444
box 5748 19444 5948 19520
use cut_M2M4_2x1 
transform 1 0 5748 0 1 20404
box 5748 20404 5948 20480
use cut_M2M4_2x1 
transform 1 0 5748 0 1 21364
box 5748 21364 5948 21440
use cut_M2M4_2x1 
transform 1 0 5748 0 1 22324
box 5748 22324 5948 22400
use cut_M2M4_2x1 
transform 1 0 5748 0 1 23284
box 5748 23284 5948 23360
use cut_M2M4_2x1 
transform 1 0 5748 0 1 24244
box 5748 24244 5948 24320
use cut_M2M4_2x1 
transform 1 0 5748 0 1 25204
box 5748 25204 5948 25280
use cut_M2M4_2x1 
transform 1 0 5748 0 1 26164
box 5748 26164 5948 26240
use cut_M2M4_2x1 
transform 1 0 5748 0 1 27124
box 5748 27124 5948 27200
use cut_M2M4_2x1 
transform 1 0 5748 0 1 28084
box 5748 28084 5948 28160
use cut_M2M4_2x1 
transform 1 0 5748 0 1 29044
box 5748 29044 5948 29120
use cut_M2M4_2x1 
transform 1 0 5748 0 1 30004
box 5748 30004 5948 30080
use cut_M2M4_2x1 
transform 1 0 5748 0 1 30964
box 5748 30964 5948 31040
use cut_M2M4_2x1 
transform 1 0 5748 0 1 31924
box 5748 31924 5948 32000
use cut_M2M4_2x1 
transform 1 0 5748 0 1 32884
box 5748 32884 5948 32960
use cut_M2M4_2x1 
transform 1 0 5748 0 1 33844
box 5748 33844 5948 33920
use cut_M2M4_2x1 
transform 1 0 5748 0 1 34804
box 5748 34804 5948 34880
use cut_M2M4_2x1 
transform 1 0 5748 0 1 35764
box 5748 35764 5948 35840
use cut_M2M4_2x1 
transform 1 0 5748 0 1 36724
box 5748 36724 5948 36800
use cut_M2M4_2x1 
transform 1 0 5748 0 1 37684
box 5748 37684 5948 37760
use cut_M2M4_2x1 
transform 1 0 5748 0 1 38644
box 5748 38644 5948 38720
use cut_M2M4_2x1 
transform 1 0 5748 0 1 39604
box 5748 39604 5948 39680
use cut_M2M4_2x1 
transform 1 0 5748 0 1 40564
box 5748 40564 5948 40640
use cut_M2M4_2x1 
transform 1 0 5748 0 1 41524
box 5748 41524 5948 41600
use cut_M2M4_2x1 
transform 1 0 5748 0 1 42484
box 5748 42484 5948 42560
use cut_M2M4_2x1 
transform 1 0 5748 0 1 43444
box 5748 43444 5948 43520
use cut_M2M4_2x1 
transform 1 0 5748 0 1 44404
box 5748 44404 5948 44480
use cut_M2M4_2x1 
transform 1 0 5748 0 1 45364
box 5748 45364 5948 45440
use cut_M2M4_2x1 
transform 1 0 5748 0 1 46324
box 5748 46324 5948 46400
use cut_M2M4_2x1 
transform 1 0 5748 0 1 47284
box 5748 47284 5948 47360
use cut_M2M4_2x1 
transform 1 0 5748 0 1 48244
box 5748 48244 5948 48320
use cut_M2M4_2x1 
transform 1 0 5748 0 1 49204
box 5748 49204 5948 49280
use cut_M1M3_2x1 
transform 1 0 1060 0 1 4058
box 1060 4058 1260 4134
use cut_M3M4_2x1 
transform 1 0 5748 0 1 1204
box 5748 1204 5948 1280
use cut_M3M4_2x1 
transform 1 0 5748 0 1 2164
box 5748 2164 5948 2240
use cut_M3M4_2x1 
transform 1 0 5748 0 1 3124
box 5748 3124 5948 3200
use cut_M1M4_1x2 
transform 1 0 39532 0 1 0
box 39532 0 39608 200
use cut_M1M4_1x2 
transform 1 0 39532 0 1 404
box 39532 404 39608 604
use cut_M1M4_1x2 
transform 1 0 39532 0 1 1364
box 39532 1364 39608 1564
use cut_M1M4_1x2 
transform 1 0 39532 0 1 2324
box 39532 2324 39608 2524
use cut_M1M4_1x2 
transform 1 0 39532 0 1 3284
box 39532 3284 39608 3484
use cut_M1M4_1x2 
transform 1 0 39532 0 1 4244
box 39532 4244 39608 4444
use cut_M1M4_1x2 
transform 1 0 39532 0 1 5204
box 39532 5204 39608 5404
use cut_M1M4_1x2 
transform 1 0 39532 0 1 6164
box 39532 6164 39608 6364
use cut_M1M4_1x2 
transform 1 0 39532 0 1 7124
box 39532 7124 39608 7324
use cut_M1M4_1x2 
transform 1 0 39532 0 1 8084
box 39532 8084 39608 8284
use cut_M1M4_1x2 
transform 1 0 39532 0 1 9044
box 39532 9044 39608 9244
use cut_M1M4_1x2 
transform 1 0 39532 0 1 10004
box 39532 10004 39608 10204
use cut_M1M4_1x2 
transform 1 0 39532 0 1 10964
box 39532 10964 39608 11164
use cut_M1M4_1x2 
transform 1 0 39532 0 1 11924
box 39532 11924 39608 12124
use cut_M1M4_1x2 
transform 1 0 39532 0 1 12884
box 39532 12884 39608 13084
use cut_M1M4_1x2 
transform 1 0 39532 0 1 13844
box 39532 13844 39608 14044
use cut_M1M4_1x2 
transform 1 0 39532 0 1 14804
box 39532 14804 39608 15004
use cut_M1M4_1x2 
transform 1 0 39532 0 1 15764
box 39532 15764 39608 15964
use cut_M1M4_1x2 
transform 1 0 39532 0 1 16724
box 39532 16724 39608 16924
use cut_M1M4_1x2 
transform 1 0 39532 0 1 17684
box 39532 17684 39608 17884
use cut_M1M4_1x2 
transform 1 0 39532 0 1 18644
box 39532 18644 39608 18844
use cut_M1M4_1x2 
transform 1 0 39532 0 1 19604
box 39532 19604 39608 19804
use cut_M1M4_1x2 
transform 1 0 39532 0 1 20564
box 39532 20564 39608 20764
use cut_M1M4_1x2 
transform 1 0 39532 0 1 21524
box 39532 21524 39608 21724
use cut_M1M4_1x2 
transform 1 0 39532 0 1 22484
box 39532 22484 39608 22684
use cut_M1M4_1x2 
transform 1 0 39532 0 1 23444
box 39532 23444 39608 23644
use cut_M1M4_1x2 
transform 1 0 39532 0 1 24404
box 39532 24404 39608 24604
use cut_M1M4_1x2 
transform 1 0 39532 0 1 25364
box 39532 25364 39608 25564
use cut_M1M4_1x2 
transform 1 0 39532 0 1 26324
box 39532 26324 39608 26524
use cut_M1M4_1x2 
transform 1 0 39532 0 1 27284
box 39532 27284 39608 27484
use cut_M1M4_1x2 
transform 1 0 39532 0 1 28244
box 39532 28244 39608 28444
use cut_M1M4_1x2 
transform 1 0 39532 0 1 29204
box 39532 29204 39608 29404
use cut_M1M4_1x2 
transform 1 0 39532 0 1 30164
box 39532 30164 39608 30364
use cut_M1M4_1x2 
transform 1 0 39532 0 1 31124
box 39532 31124 39608 31324
use cut_M1M4_1x2 
transform 1 0 39532 0 1 32084
box 39532 32084 39608 32284
use cut_M1M4_1x2 
transform 1 0 39532 0 1 33044
box 39532 33044 39608 33244
use cut_M1M4_1x2 
transform 1 0 39532 0 1 34004
box 39532 34004 39608 34204
use cut_M1M4_1x2 
transform 1 0 39532 0 1 34964
box 39532 34964 39608 35164
use cut_M1M4_1x2 
transform 1 0 39532 0 1 35924
box 39532 35924 39608 36124
use cut_M1M4_1x2 
transform 1 0 39532 0 1 36884
box 39532 36884 39608 37084
use cut_M1M4_1x2 
transform 1 0 39532 0 1 37844
box 39532 37844 39608 38044
use cut_M1M4_1x2 
transform 1 0 39532 0 1 38804
box 39532 38804 39608 39004
use cut_M1M4_1x2 
transform 1 0 39532 0 1 39764
box 39532 39764 39608 39964
use cut_M1M4_1x2 
transform 1 0 39532 0 1 40724
box 39532 40724 39608 40924
use cut_M1M4_1x2 
transform 1 0 39532 0 1 41684
box 39532 41684 39608 41884
use cut_M1M4_1x2 
transform 1 0 39532 0 1 42644
box 39532 42644 39608 42844
use cut_M1M4_1x2 
transform 1 0 39532 0 1 43604
box 39532 43604 39608 43804
use cut_M1M4_1x2 
transform 1 0 39532 0 1 44564
box 39532 44564 39608 44764
use cut_M1M4_1x2 
transform 1 0 39532 0 1 45524
box 39532 45524 39608 45724
use cut_M1M4_1x2 
transform 1 0 39532 0 1 46484
box 39532 46484 39608 46684
use cut_M1M4_1x2 
transform 1 0 39532 0 1 47444
box 39532 47444 39608 47644
use cut_M1M4_1x2 
transform 1 0 39532 0 1 48404
box 39532 48404 39608 48604
<< labels >>
flabel locali s 39532 0 39832 49848 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 4516 21706 5092 21926 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew
flabel locali s 1060 4058 1636 4278 0 FreeSans 400 0 0 0 VLPF
port 3 nsew
<< end >>
