magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 640
<< locali >>
rect 400 450 568 510
rect 568 50 800 110
rect 568 50 628 510
rect 800 50 968 110
rect 968 50 1520 110
rect 968 50 1028 110
rect 800 530 968 590
rect 968 530 1520 590
rect 968 530 1028 590
<< poly >>
rect 280 142 2040 178
rect 280 462 2040 498
<< m3 >>
rect 1400 0 1600 640
rect 680 0 880 640
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use cut_M1M4_2x1 
transform 1 0 1400 0 1 210
box 1400 210 1600 278
use cut_M1M4_2x1 
transform 1 0 1400 0 1 370
box 1400 370 1600 438
use cut_M1M4_2x1 
transform 1 0 680 0 1 210
box 680 210 880 278
use cut_M1M4_2x1 
transform 1 0 680 0 1 370
box 680 370 880 438
<< labels >>
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 680 530 920 590 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel locali s 2200 120 2440 200 0 FreeSans 400 0 0 0 BULKP
port 3 nsew
flabel locali s -120 120 120 200 0 FreeSans 400 0 0 0 BULKN
port 4 nsew
flabel m3 s 1400 0 1600 640 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 680 0 880 640 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
