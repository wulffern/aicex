magic
tech sky130A
magscale 1 2
timestamp 1659285988
<< checkpaint >>
rect 0 0 200 200
<< locali >>
rect 0 0 184 184
<< viali >>
rect 12 12 68 68
rect 12 116 68 172
rect 116 12 172 68
rect 116 116 172 172
<< m1 >>
rect 0 0 184 184
<< v1 >>
rect 12 12 68 68
rect 12 116 68 172
rect 116 12 172 68
rect 116 116 172 172
<< m2 >>
rect 0 0 200 200
<< v2 >>
rect 12 12 76 76
rect 12 124 76 188
rect 124 12 188 76
rect 124 124 188 188
<< m3 >>
rect 0 0 200 200
<< labels >>
<< end >>
