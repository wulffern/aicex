magic
tech sky130A
magscale 1 2
timestamp 1661983200
<< checkpaint >>
rect 0 0 4752 2860
<< ppolyres >>
rect 360 -110 504 110
rect 792 -110 936 110
rect 1224 -110 1368 110
rect 1656 -110 1800 110
rect 2088 -110 2232 110
rect 2520 -110 2664 110
rect 2952 -110 3096 110
rect 3384 -110 3528 110
rect 3816 -110 3960 110
rect 4248 -110 4392 110
rect 360 110 504 330
rect 792 110 936 330
rect 1224 110 1368 330
rect 1656 110 1800 330
rect 2088 110 2232 330
rect 2520 110 2664 330
rect 2952 110 3096 330
rect 3384 110 3528 330
rect 3816 110 3960 330
rect 4248 110 4392 330
rect 360 330 504 550
rect 792 330 936 550
rect 1224 330 1368 550
rect 1656 330 1800 550
rect 2088 330 2232 550
rect 2520 330 2664 550
rect 2952 330 3096 550
rect 3384 330 3528 550
rect 3816 330 3960 550
rect 4248 330 4392 550
rect 360 550 504 770
rect 792 550 936 770
rect 1224 550 1368 770
rect 1656 550 1800 770
rect 2088 550 2232 770
rect 2520 550 2664 770
rect 2952 550 3096 770
rect 3384 550 3528 770
rect 3816 550 3960 770
rect 4248 550 4392 770
rect 360 770 504 990
rect 792 770 936 990
rect 1224 770 1368 990
rect 1656 770 1800 990
rect 2088 770 2232 990
rect 2520 770 2664 990
rect 2952 770 3096 990
rect 3384 770 3528 990
rect 3816 770 3960 990
rect 4248 770 4392 990
rect 360 990 504 1210
rect 792 990 936 1210
rect 1224 990 1368 1210
rect 1656 990 1800 1210
rect 2088 990 2232 1210
rect 2520 990 2664 1210
rect 2952 990 3096 1210
rect 3384 990 3528 1210
rect 3816 990 3960 1210
rect 4248 990 4392 1210
rect 360 1210 504 1430
rect 792 1210 936 1430
rect 1224 1210 1368 1430
rect 1656 1210 1800 1430
rect 2088 1210 2232 1430
rect 2520 1210 2664 1430
rect 2952 1210 3096 1430
rect 3384 1210 3528 1430
rect 3816 1210 3960 1430
rect 4248 1210 4392 1430
rect 360 1430 504 1650
rect 792 1430 936 1650
rect 1224 1430 1368 1650
rect 1656 1430 1800 1650
rect 2088 1430 2232 1650
rect 2520 1430 2664 1650
rect 2952 1430 3096 1650
rect 3384 1430 3528 1650
rect 3816 1430 3960 1650
rect 4248 1430 4392 1650
rect 360 1650 504 1870
rect 792 1650 936 1870
rect 1224 1650 1368 1870
rect 1656 1650 1800 1870
rect 2088 1650 2232 1870
rect 2520 1650 2664 1870
rect 2952 1650 3096 1870
rect 3384 1650 3528 1870
rect 3816 1650 3960 1870
rect 4248 1650 4392 1870
rect 360 1870 504 2090
rect 792 1870 936 2090
rect 1224 1870 1368 2090
rect 1656 1870 1800 2090
rect 2088 1870 2232 2090
rect 2520 1870 2664 2090
rect 2952 1870 3096 2090
rect 3384 1870 3528 2090
rect 3816 1870 3960 2090
rect 4248 1870 4392 2090
rect 360 2090 504 2310
rect 792 2090 936 2310
rect 1224 2090 1368 2310
rect 1656 2090 1800 2310
rect 2088 2090 2232 2310
rect 2520 2090 2664 2310
rect 2952 2090 3096 2310
rect 3384 2090 3528 2310
rect 3816 2090 3960 2310
rect 4248 2090 4392 2310
rect 360 2310 504 2530
rect 792 2310 936 2530
rect 1224 2310 1368 2530
rect 1656 2310 1800 2530
rect 2088 2310 2232 2530
rect 2520 2310 2664 2530
rect 2952 2310 3096 2530
rect 3384 2310 3528 2530
rect 3816 2310 3960 2530
rect 4248 2310 4392 2530
<< poly >>
rect -72 -110 72 110
rect 4680 -110 4824 110
rect -72 110 72 330
rect 4680 110 4824 330
rect -72 330 72 550
rect 4680 330 4824 550
rect -72 550 72 770
rect 4680 550 4824 770
rect -72 770 72 990
rect 4680 770 4824 990
rect -72 990 72 1210
rect 4680 990 4824 1210
rect -72 1210 72 1430
rect 4680 1210 4824 1430
rect -72 1430 72 1650
rect 4680 1430 4824 1650
rect -72 1650 72 1870
rect 4680 1650 4824 1870
rect -72 1870 72 2090
rect 4680 1870 4824 2090
rect -72 2090 72 2310
rect 4680 2090 4824 2310
rect -72 2310 72 2530
rect 4680 2310 4824 2530
<< xpolycontact >>
rect 360 -110 504 110
rect 792 -110 936 110
rect 1224 -110 1368 110
rect 1656 -110 1800 110
rect 2088 -110 2232 110
rect 2520 -110 2664 110
rect 2952 -110 3096 110
rect 3384 -110 3528 110
rect 3816 -110 3960 110
rect 4248 -110 4392 110
rect 360 110 504 330
rect 792 110 936 330
rect 1224 110 1368 330
rect 1656 110 1800 330
rect 2088 110 2232 330
rect 2520 110 2664 330
rect 2952 110 3096 330
rect 3384 110 3528 330
rect 3816 110 3960 330
rect 4248 110 4392 330
rect 360 2090 504 2310
rect 792 2090 936 2310
rect 1224 2090 1368 2310
rect 1656 2090 1800 2310
rect 2088 2090 2232 2310
rect 2520 2090 2664 2310
rect 2952 2090 3096 2310
rect 3384 2090 3528 2310
rect 3816 2090 3960 2310
rect 4248 2090 4392 2310
rect 360 2310 504 2530
rect 792 2310 936 2530
rect 1224 2310 1368 2530
rect 1656 2310 1800 2530
rect 2088 2310 2232 2530
rect 2520 2310 2664 2530
rect 2952 2310 3096 2530
rect 3384 2310 3528 2530
rect 3816 2310 3960 2530
rect 4248 2310 4392 2530
<< locali >>
rect 360 -110 936 110
rect 1224 -110 1800 110
rect 2088 -110 2664 110
rect 2952 -110 3528 110
rect 3816 -110 4392 110
rect 360 110 936 330
rect 1224 110 1800 330
rect 2088 110 2664 330
rect 2952 110 3528 330
rect 3816 110 4392 330
rect 360 2090 504 2310
rect 792 2090 936 2310
rect 1224 2090 1368 2310
rect 1656 2090 1800 2310
rect 2088 2090 2232 2310
rect 2520 2090 2664 2310
rect 2952 2090 3096 2310
rect 3384 2090 3528 2310
rect 3816 2090 3960 2310
rect 4248 2090 4392 2310
rect 360 2310 504 2530
rect 792 2310 936 2530
rect 1224 2310 1368 2530
rect 1656 2310 1800 2530
rect 2088 2310 2232 2530
rect 2520 2310 2664 2530
rect 2952 2310 3096 2530
rect 3384 2310 3528 2530
rect 3816 2310 3960 2530
rect 4248 2310 4392 2530
rect 360 2530 504 2750
rect 792 2530 936 2750
rect 1224 2530 1368 2750
rect 1656 2530 1800 2750
rect 2088 2530 2232 2750
rect 2520 2530 2664 2750
rect 2952 2530 3096 2750
rect 3384 2530 3528 2750
rect 3816 2530 3960 2750
rect 4248 2530 4392 2750
rect -72 2750 504 2970
rect -72 2750 504 2970
rect 792 2750 1368 2970
rect 1656 2750 2232 2970
rect 2520 2750 3096 2970
rect 3384 2750 3960 2970
rect 4248 2750 4824 2970
rect 4248 2750 4824 2970
<< pwell >>
rect -72 -110 4824 2970
<< labels >>
flabel locali s -72 2750 504 2970 0 FreeSans 400 0 0 0 N
port 1 nsew
flabel locali s 4248 2750 4824 2970 0 FreeSans 400 0 0 0 P
port 2 nsew
<< end >>
