magic
tech sky130A
magscale 1 2
timestamp 1658582973
<< checkpaint >>
rect 0 0 200 76
<< m3 >>
rect 0 0 200 76
<< m4 >>
rect 0 0 200 76
<< v3 >>
rect 12 6 188 70
<< labels >>
<< end >>
