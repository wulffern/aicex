magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 11280 960
<< m1 >>
rect 120 -40 11240 40
rect 11160 40 11240 120
rect 120 120 11080 200
rect 11160 120 11240 200
rect 120 200 200 280
rect 11160 200 11240 280
rect 120 280 200 360
rect 280 280 11240 360
rect 120 360 200 440
rect 11160 360 11240 440
rect 120 440 11080 520
rect 11160 440 11240 520
rect 120 520 200 600
rect 11160 520 11240 600
rect 120 600 200 680
rect 280 600 11240 680
rect 120 680 200 760
rect 120 760 11240 840
<< m2 >>
rect 120 -40 11240 40
rect 11160 40 11240 120
rect 120 120 11080 200
rect 11160 120 11240 200
rect 120 200 200 280
rect 11160 200 11240 280
rect 120 280 200 360
rect 280 280 11240 360
rect 120 360 200 440
rect 11160 360 11240 440
rect 120 440 11080 520
rect 11160 440 11240 520
rect 120 520 200 600
rect 11160 520 11240 600
rect 120 600 200 680
rect 280 600 11240 680
rect 120 680 200 760
rect 120 760 11240 840
<< locali >>
rect 120 -40 11240 40
rect 11160 40 11240 120
rect 120 120 11080 200
rect 11160 120 11240 200
rect 120 200 200 280
rect 11160 200 11240 280
rect 120 280 200 360
rect 280 280 11240 360
rect 120 360 200 440
rect 11160 360 11240 440
rect 120 440 11080 520
rect 11160 440 11240 520
rect 120 520 200 600
rect 11160 520 11240 600
rect 120 600 200 680
rect 280 600 11240 680
rect 120 680 200 760
rect 120 760 11240 840
<< v1 >>
rect 10840 -32 10919 -24
rect 10840 -24 10919 -16
rect 10840 -16 10919 -8
rect 10840 -8 10919 0
rect 10840 0 10919 8
rect 10840 8 10919 16
rect 10840 16 10919 24
rect 10840 24 10919 32
rect 10920 -32 10999 -24
rect 10920 -24 10999 -16
rect 10920 -16 10999 -8
rect 10920 -8 10999 0
rect 10920 0 10999 8
rect 10920 8 10999 16
rect 10920 16 10999 24
rect 10920 24 10999 32
rect 11000 -32 11079 -24
rect 11000 -24 11079 -16
rect 11000 -16 11079 -8
rect 11000 -8 11079 0
rect 11000 0 11079 8
rect 11000 8 11079 16
rect 11000 16 11079 24
rect 11000 24 11079 32
rect 360 128 439 136
rect 360 136 439 144
rect 360 144 439 152
rect 360 152 439 160
rect 360 160 439 168
rect 360 168 439 176
rect 360 176 439 184
rect 360 184 439 192
rect 440 128 519 136
rect 440 136 519 144
rect 440 144 519 152
rect 440 152 519 160
rect 440 160 519 168
rect 440 168 519 176
rect 440 176 519 184
rect 440 184 519 192
rect 520 128 599 136
rect 520 136 599 144
rect 520 144 599 152
rect 520 152 599 160
rect 520 160 599 168
rect 520 168 599 176
rect 520 176 599 184
rect 520 184 599 192
rect 10840 288 10919 296
rect 10840 296 10919 304
rect 10840 304 10919 312
rect 10840 312 10919 320
rect 10840 320 10919 328
rect 10840 328 10919 336
rect 10840 336 10919 344
rect 10840 344 10919 352
rect 10920 288 10999 296
rect 10920 296 10999 304
rect 10920 304 10999 312
rect 10920 312 10999 320
rect 10920 320 10999 328
rect 10920 328 10999 336
rect 10920 336 10999 344
rect 10920 344 10999 352
rect 11000 288 11079 296
rect 11000 296 11079 304
rect 11000 304 11079 312
rect 11000 312 11079 320
rect 11000 320 11079 328
rect 11000 328 11079 336
rect 11000 336 11079 344
rect 11000 344 11079 352
rect 360 448 439 456
rect 360 456 439 464
rect 360 464 439 472
rect 360 472 439 480
rect 360 480 439 488
rect 360 488 439 496
rect 360 496 439 504
rect 360 504 439 512
rect 440 448 519 456
rect 440 456 519 464
rect 440 464 519 472
rect 440 472 519 480
rect 440 480 519 488
rect 440 488 519 496
rect 440 496 519 504
rect 440 504 519 512
rect 520 448 599 456
rect 520 456 599 464
rect 520 464 599 472
rect 520 472 599 480
rect 520 480 599 488
rect 520 488 599 496
rect 520 496 599 504
rect 520 504 599 512
rect 10840 608 10919 616
rect 10840 616 10919 624
rect 10840 624 10919 632
rect 10840 632 10919 640
rect 10840 640 10919 648
rect 10840 648 10919 656
rect 10840 656 10919 664
rect 10840 664 10919 672
rect 10920 608 10999 616
rect 10920 616 10999 624
rect 10920 624 10999 632
rect 10920 632 10999 640
rect 10920 640 10999 648
rect 10920 648 10999 656
rect 10920 656 10999 664
rect 10920 664 10999 672
rect 11000 608 11079 616
rect 11000 616 11079 624
rect 11000 624 11079 632
rect 11000 632 11079 640
rect 11000 640 11079 648
rect 11000 648 11079 656
rect 11000 656 11079 664
rect 11000 664 11079 672
rect 360 768 439 776
rect 360 776 439 784
rect 360 784 439 792
rect 360 792 439 800
rect 360 800 439 808
rect 360 808 439 816
rect 360 816 439 824
rect 360 824 439 832
rect 440 768 519 776
rect 440 776 519 784
rect 440 784 519 792
rect 440 792 519 800
rect 440 800 519 808
rect 440 808 519 816
rect 440 816 519 824
rect 440 824 519 832
rect 520 768 599 776
rect 520 776 599 784
rect 520 784 599 792
rect 520 792 599 800
rect 520 800 599 808
rect 520 808 599 816
rect 520 816 599 824
rect 520 824 599 832
<< v2 >>
rect 10840 -32 10919 -24
rect 10840 -24 10919 -16
rect 10840 -16 10919 -8
rect 10840 -8 10919 0
rect 10840 0 10919 8
rect 10840 8 10919 16
rect 10840 16 10919 24
rect 10840 24 10919 32
rect 10920 -32 10999 -24
rect 10920 -24 10999 -16
rect 10920 -16 10999 -8
rect 10920 -8 10999 0
rect 10920 0 10999 8
rect 10920 8 10999 16
rect 10920 16 10999 24
rect 10920 24 10999 32
rect 11000 -32 11079 -24
rect 11000 -24 11079 -16
rect 11000 -16 11079 -8
rect 11000 -8 11079 0
rect 11000 0 11079 8
rect 11000 8 11079 16
rect 11000 16 11079 24
rect 11000 24 11079 32
rect 360 128 439 136
rect 360 136 439 144
rect 360 144 439 152
rect 360 152 439 160
rect 360 160 439 168
rect 360 168 439 176
rect 360 176 439 184
rect 360 184 439 192
rect 440 128 519 136
rect 440 136 519 144
rect 440 144 519 152
rect 440 152 519 160
rect 440 160 519 168
rect 440 168 519 176
rect 440 176 519 184
rect 440 184 519 192
rect 520 128 599 136
rect 520 136 599 144
rect 520 144 599 152
rect 520 152 599 160
rect 520 160 599 168
rect 520 168 599 176
rect 520 176 599 184
rect 520 184 599 192
rect 10840 288 10919 296
rect 10840 296 10919 304
rect 10840 304 10919 312
rect 10840 312 10919 320
rect 10840 320 10919 328
rect 10840 328 10919 336
rect 10840 336 10919 344
rect 10840 344 10919 352
rect 10920 288 10999 296
rect 10920 296 10999 304
rect 10920 304 10999 312
rect 10920 312 10999 320
rect 10920 320 10999 328
rect 10920 328 10999 336
rect 10920 336 10999 344
rect 10920 344 10999 352
rect 11000 288 11079 296
rect 11000 296 11079 304
rect 11000 304 11079 312
rect 11000 312 11079 320
rect 11000 320 11079 328
rect 11000 328 11079 336
rect 11000 336 11079 344
rect 11000 344 11079 352
rect 360 448 439 456
rect 360 456 439 464
rect 360 464 439 472
rect 360 472 439 480
rect 360 480 439 488
rect 360 488 439 496
rect 360 496 439 504
rect 360 504 439 512
rect 440 448 519 456
rect 440 456 519 464
rect 440 464 519 472
rect 440 472 519 480
rect 440 480 519 488
rect 440 488 519 496
rect 440 496 519 504
rect 440 504 519 512
rect 520 448 599 456
rect 520 456 599 464
rect 520 464 599 472
rect 520 472 599 480
rect 520 480 599 488
rect 520 488 599 496
rect 520 496 599 504
rect 520 504 599 512
rect 10840 608 10919 616
rect 10840 616 10919 624
rect 10840 624 10919 632
rect 10840 632 10919 640
rect 10840 640 10919 648
rect 10840 648 10919 656
rect 10840 656 10919 664
rect 10840 664 10919 672
rect 10920 608 10999 616
rect 10920 616 10999 624
rect 10920 624 10999 632
rect 10920 632 10999 640
rect 10920 640 10999 648
rect 10920 648 10999 656
rect 10920 656 10999 664
rect 10920 664 10999 672
rect 11000 608 11079 616
rect 11000 616 11079 624
rect 11000 624 11079 632
rect 11000 632 11079 640
rect 11000 640 11079 648
rect 11000 648 11079 656
rect 11000 656 11079 664
rect 11000 664 11079 672
rect 360 768 439 776
rect 360 776 439 784
rect 360 784 439 792
rect 360 792 439 800
rect 360 800 439 808
rect 360 808 439 816
rect 360 816 439 824
rect 360 824 439 832
rect 440 768 519 776
rect 440 776 519 784
rect 440 784 519 792
rect 440 792 519 800
rect 440 800 519 808
rect 440 808 519 816
rect 440 816 519 824
rect 440 824 519 832
rect 520 768 599 776
rect 520 776 599 784
rect 520 784 599 792
rect 520 792 599 800
rect 520 800 599 808
rect 520 808 599 816
rect 520 816 599 824
rect 520 824 599 832
<< viali >>
rect 10840 -32 10919 -24
rect 10840 -24 10919 -16
rect 10840 -16 10919 -8
rect 10840 -8 10919 0
rect 10840 0 10919 8
rect 10840 8 10919 16
rect 10840 16 10919 24
rect 10840 24 10919 32
rect 10920 -32 10999 -24
rect 10920 -24 10999 -16
rect 10920 -16 10999 -8
rect 10920 -8 10999 0
rect 10920 0 10999 8
rect 10920 8 10999 16
rect 10920 16 10999 24
rect 10920 24 10999 32
rect 11000 -32 11079 -24
rect 11000 -24 11079 -16
rect 11000 -16 11079 -8
rect 11000 -8 11079 0
rect 11000 0 11079 8
rect 11000 8 11079 16
rect 11000 16 11079 24
rect 11000 24 11079 32
rect 360 128 439 136
rect 360 136 439 144
rect 360 144 439 152
rect 360 152 439 160
rect 360 160 439 168
rect 360 168 439 176
rect 360 176 439 184
rect 360 184 439 192
rect 440 128 519 136
rect 440 136 519 144
rect 440 144 519 152
rect 440 152 519 160
rect 440 160 519 168
rect 440 168 519 176
rect 440 176 519 184
rect 440 184 519 192
rect 520 128 599 136
rect 520 136 599 144
rect 520 144 599 152
rect 520 152 599 160
rect 520 160 599 168
rect 520 168 599 176
rect 520 176 599 184
rect 520 184 599 192
rect 10840 288 10919 296
rect 10840 296 10919 304
rect 10840 304 10919 312
rect 10840 312 10919 320
rect 10840 320 10919 328
rect 10840 328 10919 336
rect 10840 336 10919 344
rect 10840 344 10919 352
rect 10920 288 10999 296
rect 10920 296 10999 304
rect 10920 304 10999 312
rect 10920 312 10999 320
rect 10920 320 10999 328
rect 10920 328 10999 336
rect 10920 336 10999 344
rect 10920 344 10999 352
rect 11000 288 11079 296
rect 11000 296 11079 304
rect 11000 304 11079 312
rect 11000 312 11079 320
rect 11000 320 11079 328
rect 11000 328 11079 336
rect 11000 336 11079 344
rect 11000 344 11079 352
rect 360 448 439 456
rect 360 456 439 464
rect 360 464 439 472
rect 360 472 439 480
rect 360 480 439 488
rect 360 488 439 496
rect 360 496 439 504
rect 360 504 439 512
rect 440 448 519 456
rect 440 456 519 464
rect 440 464 519 472
rect 440 472 519 480
rect 440 480 519 488
rect 440 488 519 496
rect 440 496 519 504
rect 440 504 519 512
rect 520 448 599 456
rect 520 456 599 464
rect 520 464 599 472
rect 520 472 599 480
rect 520 480 599 488
rect 520 488 599 496
rect 520 496 599 504
rect 520 504 599 512
rect 10840 608 10919 616
rect 10840 616 10919 624
rect 10840 624 10919 632
rect 10840 632 10919 640
rect 10840 640 10919 648
rect 10840 648 10919 656
rect 10840 656 10919 664
rect 10840 664 10919 672
rect 10920 608 10999 616
rect 10920 616 10999 624
rect 10920 624 10999 632
rect 10920 632 10999 640
rect 10920 640 10999 648
rect 10920 648 10999 656
rect 10920 656 10999 664
rect 10920 664 10999 672
rect 11000 608 11079 616
rect 11000 616 11079 624
rect 11000 624 11079 632
rect 11000 632 11079 640
rect 11000 640 11079 648
rect 11000 648 11079 656
rect 11000 656 11079 664
rect 11000 664 11079 672
rect 360 768 439 776
rect 360 776 439 784
rect 360 784 439 792
rect 360 792 439 800
rect 360 800 439 808
rect 360 808 439 816
rect 360 816 439 824
rect 360 824 439 832
rect 440 768 519 776
rect 440 776 519 784
rect 440 784 519 792
rect 440 792 519 800
rect 440 800 519 808
rect 440 808 519 816
rect 440 816 519 824
rect 440 824 519 832
rect 520 768 599 776
rect 520 776 599 784
rect 520 784 599 792
rect 520 792 599 800
rect 520 800 599 808
rect 520 808 599 816
rect 520 816 599 824
rect 520 824 599 832
<< m3 >>
rect 120 -40 11240 40
rect 11160 40 11240 120
rect 120 120 10840 200
rect 10920 120 11080 200
rect 11160 120 11240 200
rect 120 200 200 280
rect 11160 200 11240 280
rect 120 280 200 360
rect 280 280 360 360
rect 440 280 11240 360
rect 120 360 200 440
rect 11160 360 11240 440
rect 120 440 11080 520
rect 11160 440 11240 520
rect 120 520 200 600
rect 11160 520 11240 600
rect 120 600 200 680
rect 280 600 11240 680
rect 120 680 200 760
rect 120 760 11240 840
<< rm3 >>
rect 10840 120 10920 200
rect 360 280 440 360
<< labels >>
flabel m3 s 120 -40 11240 40 0 FreeSans 400 0 0 0 B
port 1 nsew
flabel m3 s 120 760 11240 840 0 FreeSans 400 0 0 0 A
port 2 nsew
<< end >>
