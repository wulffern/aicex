magic
tech sky130A
magscale 1 2
timestamp 1658600916
<< checkpaint >>
rect 112 0 11844 12540
<< m1 >>
rect 2100 4820 2160 12480
rect 2100 4820 2160 12480
rect 1920 140 1980 12480
rect 1920 140 1980 12480
rect 1740 9500 1800 12480
rect 1740 9500 1800 12480
rect 1560 1700 1620 12480
rect 1560 1700 1620 12480
rect 1380 3488 1440 12480
rect 1380 3488 1440 12480
rect 1200 8168 1260 12480
rect 1200 8168 1260 12480
rect 1020 7940 1080 12480
rect 1020 7940 1080 12480
rect 840 8624 900 12480
rect 840 8624 900 12480
rect 660 3944 720 12480
rect 660 3944 720 12480
rect 480 4172 540 12480
rect 480 4172 540 12480
rect 300 3716 360 12480
rect 300 3716 360 12480
rect 120 4400 180 12480
rect 120 4400 180 12480
rect 2668 0 11768 76
<< m2 >>
rect 2160 4882 2340 4958
rect 2160 6022 2340 6098
rect 2160 5338 2340 5414
rect 2160 5794 2340 5870
rect 2160 5566 2340 5642
rect 2160 5110 2340 5186
rect 2160 4882 2340 4958
rect 2160 6022 2340 6098
rect 2160 5338 2340 5414
rect 2160 5794 2340 5870
rect 2160 5566 2340 5642
rect 2160 5110 2340 5186
rect 2160 4882 2340 4958
rect 2160 6022 2340 6098
rect 2160 5338 2340 5414
rect 2160 5794 2340 5870
rect 2160 5566 2340 5642
rect 2160 5110 2340 5186
rect 2160 4882 2340 4958
rect 2160 6022 2340 6098
rect 2160 5338 2340 5414
rect 2160 5794 2340 5870
rect 2160 5566 2340 5642
rect 2160 5110 2340 5186
rect 2160 4882 2340 4958
rect 2160 6022 2340 6098
rect 2160 5338 2340 5414
rect 2160 5794 2340 5870
rect 2160 5566 2340 5642
rect 2160 5110 2340 5186
rect 2160 4882 2340 4958
rect 2160 6022 2340 6098
rect 2160 5338 2340 5414
rect 2160 5794 2340 5870
rect 2160 5566 2340 5642
rect 2160 5110 2340 5186
rect 2160 11122 2340 11198
rect 2160 12262 2340 12338
rect 2160 11578 2340 11654
rect 2160 12034 2340 12110
rect 2160 11806 2340 11882
rect 2160 11350 2340 11426
rect 2160 11122 2340 11198
rect 2160 12262 2340 12338
rect 2160 11578 2340 11654
rect 2160 12034 2340 12110
rect 2160 11806 2340 11882
rect 2160 11350 2340 11426
rect 2160 11122 2340 11198
rect 2160 12262 2340 12338
rect 2160 11578 2340 11654
rect 2160 12034 2340 12110
rect 2160 11806 2340 11882
rect 2160 11350 2340 11426
rect 2160 11122 2340 11198
rect 2160 12262 2340 12338
rect 2160 11578 2340 11654
rect 2160 12034 2340 12110
rect 2160 11806 2340 11882
rect 2160 11350 2340 11426
rect 2160 11122 2340 11198
rect 2160 12262 2340 12338
rect 2160 11578 2340 11654
rect 2160 12034 2340 12110
rect 2160 11806 2340 11882
rect 2160 11350 2340 11426
rect 2160 11122 2340 11198
rect 2160 12262 2340 12338
rect 2160 11578 2340 11654
rect 2160 12034 2340 12110
rect 2160 11806 2340 11882
rect 2160 11350 2340 11426
rect 1980 202 2340 278
rect 1980 1342 2340 1418
rect 1980 658 2340 734
rect 1980 1114 2340 1190
rect 1980 886 2340 962
rect 1980 430 2340 506
rect 1980 202 2340 278
rect 1980 1342 2340 1418
rect 1980 658 2340 734
rect 1980 1114 2340 1190
rect 1980 886 2340 962
rect 1980 430 2340 506
rect 1980 202 2340 278
rect 1980 1342 2340 1418
rect 1980 658 2340 734
rect 1980 1114 2340 1190
rect 1980 886 2340 962
rect 1980 430 2340 506
rect 1980 202 2340 278
rect 1980 1342 2340 1418
rect 1980 658 2340 734
rect 1980 1114 2340 1190
rect 1980 886 2340 962
rect 1980 430 2340 506
rect 1980 202 2340 278
rect 1980 1342 2340 1418
rect 1980 658 2340 734
rect 1980 1114 2340 1190
rect 1980 886 2340 962
rect 1980 430 2340 506
rect 1980 202 2340 278
rect 1980 1342 2340 1418
rect 1980 658 2340 734
rect 1980 1114 2340 1190
rect 1980 886 2340 962
rect 1980 430 2340 506
rect 1980 6442 2340 6518
rect 1980 7582 2340 7658
rect 1980 6898 2340 6974
rect 1980 7354 2340 7430
rect 1980 7126 2340 7202
rect 1980 6670 2340 6746
rect 1980 6442 2340 6518
rect 1980 7582 2340 7658
rect 1980 6898 2340 6974
rect 1980 7354 2340 7430
rect 1980 7126 2340 7202
rect 1980 6670 2340 6746
rect 1980 6442 2340 6518
rect 1980 7582 2340 7658
rect 1980 6898 2340 6974
rect 1980 7354 2340 7430
rect 1980 7126 2340 7202
rect 1980 6670 2340 6746
rect 1980 6442 2340 6518
rect 1980 7582 2340 7658
rect 1980 6898 2340 6974
rect 1980 7354 2340 7430
rect 1980 7126 2340 7202
rect 1980 6670 2340 6746
rect 1980 6442 2340 6518
rect 1980 7582 2340 7658
rect 1980 6898 2340 6974
rect 1980 7354 2340 7430
rect 1980 7126 2340 7202
rect 1980 6670 2340 6746
rect 1980 6442 2340 6518
rect 1980 7582 2340 7658
rect 1980 6898 2340 6974
rect 1980 7354 2340 7430
rect 1980 7126 2340 7202
rect 1980 6670 2340 6746
rect 1800 9562 2340 9638
rect 1800 10702 2340 10778
rect 1800 10018 2340 10094
rect 1800 10474 2340 10550
rect 1800 10246 2340 10322
rect 1800 9790 2340 9866
rect 1800 9562 2340 9638
rect 1800 10702 2340 10778
rect 1800 10018 2340 10094
rect 1800 10474 2340 10550
rect 1800 10246 2340 10322
rect 1800 9790 2340 9866
rect 1800 9562 2340 9638
rect 1800 10702 2340 10778
rect 1800 10018 2340 10094
rect 1800 10474 2340 10550
rect 1800 10246 2340 10322
rect 1800 9790 2340 9866
rect 1800 9562 2340 9638
rect 1800 10702 2340 10778
rect 1800 10018 2340 10094
rect 1800 10474 2340 10550
rect 1800 10246 2340 10322
rect 1800 9790 2340 9866
rect 1800 9562 2340 9638
rect 1800 10702 2340 10778
rect 1800 10018 2340 10094
rect 1800 10474 2340 10550
rect 1800 10246 2340 10322
rect 1800 9790 2340 9866
rect 1800 9562 2340 9638
rect 1800 10702 2340 10778
rect 1800 10018 2340 10094
rect 1800 10474 2340 10550
rect 1800 10246 2340 10322
rect 1800 9790 2340 9866
rect 1620 1762 2340 1838
rect 1620 2902 2340 2978
rect 1620 2218 2340 2294
rect 1620 2674 2340 2750
rect 1620 2446 2340 2522
rect 1620 1990 2340 2066
rect 1620 1762 2340 1838
rect 1620 2902 2340 2978
rect 1620 2218 2340 2294
rect 1620 2674 2340 2750
rect 1620 2446 2340 2522
rect 1620 1990 2340 2066
rect 1620 1762 2340 1838
rect 1620 2902 2340 2978
rect 1620 2218 2340 2294
rect 1620 2674 2340 2750
rect 1620 2446 2340 2522
rect 1620 1990 2340 2066
rect 1620 1762 2340 1838
rect 1620 2902 2340 2978
rect 1620 2218 2340 2294
rect 1620 2674 2340 2750
rect 1620 2446 2340 2522
rect 1620 1990 2340 2066
rect 1620 1762 2340 1838
rect 1620 2902 2340 2978
rect 1620 2218 2340 2294
rect 1620 2674 2340 2750
rect 1620 2446 2340 2522
rect 1620 1990 2340 2066
rect 1620 1762 2340 1838
rect 1620 2902 2340 2978
rect 1620 2218 2340 2294
rect 1620 2674 2340 2750
rect 1620 2446 2340 2522
rect 1620 1990 2340 2066
rect 1440 3550 2340 3626
rect 1260 8230 2340 8306
rect 1080 8002 2340 8078
rect 1080 9142 2340 9218
rect 1080 8458 2340 8534
rect 1080 8914 2340 8990
rect 1080 8002 2340 8078
rect 1080 9142 2340 9218
rect 1080 8458 2340 8534
rect 1080 8914 2340 8990
rect 1080 8002 2340 8078
rect 1080 9142 2340 9218
rect 1080 8458 2340 8534
rect 1080 8914 2340 8990
rect 1080 8002 2340 8078
rect 1080 9142 2340 9218
rect 1080 8458 2340 8534
rect 1080 8914 2340 8990
rect 900 8686 2340 8762
rect 720 4006 2340 4082
rect 540 4234 2340 4310
rect 360 3778 2340 3854
rect 180 4462 2340 4538
<< m3 >>
rect 2668 10920 2744 12540
use CAP32C_CV XC1
transform 1 0 2340 0 1 0
box 2340 0 11844 1560
use CAP32C_CV XC64a<0>
transform 1 0 2340 0 1 1560
box 2340 1560 11844 3120
use CAP32C_CV XC32a<0>
transform 1 0 2340 0 1 3120
box 2340 3120 11844 4680
use CAP32C_CV XC128a<1>
transform 1 0 2340 0 1 4680
box 2340 4680 11844 6240
use CAP32C_CV XC128b<2>
transform 1 0 2340 0 1 6240
box 2340 6240 11844 7800
use CAP32C_CV X16ab
transform 1 0 2340 0 1 7800
box 2340 7800 11844 9360
use CAP32C_CV XC64b<1>
transform 1 0 2340 0 1 9360
box 2340 9360 11844 10920
use CAP32C_CV XC0
transform 1 0 2340 0 1 10920
box 2340 10920 11844 12480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4882
box 2340 4882 2540 4958
use cut_M2M3_1x2 
transform 1 0 2092 0 1 4820
box 2092 4820 2168 5020
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6022
box 2340 6022 2540 6098
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5960
box 2092 5960 2168 6160
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5338
box 2340 5338 2540 5414
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5276
box 2092 5276 2168 5476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5794
box 2340 5794 2540 5870
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5732
box 2092 5732 2168 5932
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5566
box 2340 5566 2540 5642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5504
box 2092 5504 2168 5704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5110
box 2340 5110 2540 5186
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5048
box 2092 5048 2168 5248
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4882
box 2340 4882 2540 4958
use cut_M2M3_1x2 
transform 1 0 2092 0 1 4820
box 2092 4820 2168 5020
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6022
box 2340 6022 2540 6098
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5960
box 2092 5960 2168 6160
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5338
box 2340 5338 2540 5414
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5276
box 2092 5276 2168 5476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5794
box 2340 5794 2540 5870
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5732
box 2092 5732 2168 5932
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5566
box 2340 5566 2540 5642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5504
box 2092 5504 2168 5704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5110
box 2340 5110 2540 5186
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5048
box 2092 5048 2168 5248
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4882
box 2340 4882 2540 4958
use cut_M2M3_1x2 
transform 1 0 2092 0 1 4820
box 2092 4820 2168 5020
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6022
box 2340 6022 2540 6098
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5960
box 2092 5960 2168 6160
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5338
box 2340 5338 2540 5414
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5276
box 2092 5276 2168 5476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5794
box 2340 5794 2540 5870
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5732
box 2092 5732 2168 5932
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5566
box 2340 5566 2540 5642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5504
box 2092 5504 2168 5704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5110
box 2340 5110 2540 5186
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5048
box 2092 5048 2168 5248
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4882
box 2340 4882 2540 4958
use cut_M2M3_1x2 
transform 1 0 2092 0 1 4820
box 2092 4820 2168 5020
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6022
box 2340 6022 2540 6098
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5960
box 2092 5960 2168 6160
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5338
box 2340 5338 2540 5414
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5276
box 2092 5276 2168 5476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5794
box 2340 5794 2540 5870
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5732
box 2092 5732 2168 5932
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5566
box 2340 5566 2540 5642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5504
box 2092 5504 2168 5704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5110
box 2340 5110 2540 5186
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5048
box 2092 5048 2168 5248
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4882
box 2340 4882 2540 4958
use cut_M2M3_1x2 
transform 1 0 2092 0 1 4820
box 2092 4820 2168 5020
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6022
box 2340 6022 2540 6098
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5960
box 2092 5960 2168 6160
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5338
box 2340 5338 2540 5414
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5276
box 2092 5276 2168 5476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5794
box 2340 5794 2540 5870
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5732
box 2092 5732 2168 5932
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5566
box 2340 5566 2540 5642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5504
box 2092 5504 2168 5704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5110
box 2340 5110 2540 5186
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5048
box 2092 5048 2168 5248
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4882
box 2340 4882 2540 4958
use cut_M2M3_1x2 
transform 1 0 2092 0 1 4820
box 2092 4820 2168 5020
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6022
box 2340 6022 2540 6098
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5960
box 2092 5960 2168 6160
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5338
box 2340 5338 2540 5414
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5276
box 2092 5276 2168 5476
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5794
box 2340 5794 2540 5870
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5732
box 2092 5732 2168 5932
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5566
box 2340 5566 2540 5642
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5504
box 2092 5504 2168 5704
use cut_M1M3_2x1 
transform 1 0 2340 0 1 5110
box 2340 5110 2540 5186
use cut_M2M3_1x2 
transform 1 0 2092 0 1 5048
box 2092 5048 2168 5248
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11122
box 2340 11122 2540 11198
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11060
box 2092 11060 2168 11260
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12262
box 2340 12262 2540 12338
use cut_M2M3_1x2 
transform 1 0 2092 0 1 12200
box 2092 12200 2168 12400
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11578
box 2340 11578 2540 11654
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11516
box 2092 11516 2168 11716
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12034
box 2340 12034 2540 12110
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11972
box 2092 11972 2168 12172
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11806
box 2340 11806 2540 11882
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11744
box 2092 11744 2168 11944
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11350
box 2340 11350 2540 11426
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11288
box 2092 11288 2168 11488
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11122
box 2340 11122 2540 11198
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11060
box 2092 11060 2168 11260
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12262
box 2340 12262 2540 12338
use cut_M2M3_1x2 
transform 1 0 2092 0 1 12200
box 2092 12200 2168 12400
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11578
box 2340 11578 2540 11654
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11516
box 2092 11516 2168 11716
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12034
box 2340 12034 2540 12110
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11972
box 2092 11972 2168 12172
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11806
box 2340 11806 2540 11882
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11744
box 2092 11744 2168 11944
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11350
box 2340 11350 2540 11426
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11288
box 2092 11288 2168 11488
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11122
box 2340 11122 2540 11198
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11060
box 2092 11060 2168 11260
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12262
box 2340 12262 2540 12338
use cut_M2M3_1x2 
transform 1 0 2092 0 1 12200
box 2092 12200 2168 12400
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11578
box 2340 11578 2540 11654
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11516
box 2092 11516 2168 11716
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12034
box 2340 12034 2540 12110
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11972
box 2092 11972 2168 12172
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11806
box 2340 11806 2540 11882
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11744
box 2092 11744 2168 11944
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11350
box 2340 11350 2540 11426
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11288
box 2092 11288 2168 11488
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11122
box 2340 11122 2540 11198
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11060
box 2092 11060 2168 11260
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12262
box 2340 12262 2540 12338
use cut_M2M3_1x2 
transform 1 0 2092 0 1 12200
box 2092 12200 2168 12400
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11578
box 2340 11578 2540 11654
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11516
box 2092 11516 2168 11716
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12034
box 2340 12034 2540 12110
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11972
box 2092 11972 2168 12172
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11806
box 2340 11806 2540 11882
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11744
box 2092 11744 2168 11944
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11350
box 2340 11350 2540 11426
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11288
box 2092 11288 2168 11488
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11122
box 2340 11122 2540 11198
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11060
box 2092 11060 2168 11260
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12262
box 2340 12262 2540 12338
use cut_M2M3_1x2 
transform 1 0 2092 0 1 12200
box 2092 12200 2168 12400
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11578
box 2340 11578 2540 11654
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11516
box 2092 11516 2168 11716
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12034
box 2340 12034 2540 12110
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11972
box 2092 11972 2168 12172
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11806
box 2340 11806 2540 11882
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11744
box 2092 11744 2168 11944
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11350
box 2340 11350 2540 11426
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11288
box 2092 11288 2168 11488
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11122
box 2340 11122 2540 11198
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11060
box 2092 11060 2168 11260
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12262
box 2340 12262 2540 12338
use cut_M2M3_1x2 
transform 1 0 2092 0 1 12200
box 2092 12200 2168 12400
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11578
box 2340 11578 2540 11654
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11516
box 2092 11516 2168 11716
use cut_M1M3_2x1 
transform 1 0 2340 0 1 12034
box 2340 12034 2540 12110
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11972
box 2092 11972 2168 12172
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11806
box 2340 11806 2540 11882
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11744
box 2092 11744 2168 11944
use cut_M1M3_2x1 
transform 1 0 2340 0 1 11350
box 2340 11350 2540 11426
use cut_M2M3_1x2 
transform 1 0 2092 0 1 11288
box 2092 11288 2168 11488
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1342
box 2340 1342 2540 1418
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1280
box 1912 1280 1988 1480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 658
box 2340 658 2540 734
use cut_M2M3_1x2 
transform 1 0 1912 0 1 596
box 1912 596 1988 796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1114
box 2340 1114 2540 1190
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1052
box 1912 1052 1988 1252
use cut_M1M3_2x1 
transform 1 0 2340 0 1 886
box 2340 886 2540 962
use cut_M2M3_1x2 
transform 1 0 1912 0 1 824
box 1912 824 1988 1024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 430
box 2340 430 2540 506
use cut_M2M3_1x2 
transform 1 0 1912 0 1 368
box 1912 368 1988 568
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1342
box 2340 1342 2540 1418
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1280
box 1912 1280 1988 1480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 658
box 2340 658 2540 734
use cut_M2M3_1x2 
transform 1 0 1912 0 1 596
box 1912 596 1988 796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1114
box 2340 1114 2540 1190
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1052
box 1912 1052 1988 1252
use cut_M1M3_2x1 
transform 1 0 2340 0 1 886
box 2340 886 2540 962
use cut_M2M3_1x2 
transform 1 0 1912 0 1 824
box 1912 824 1988 1024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 430
box 2340 430 2540 506
use cut_M2M3_1x2 
transform 1 0 1912 0 1 368
box 1912 368 1988 568
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1342
box 2340 1342 2540 1418
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1280
box 1912 1280 1988 1480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 658
box 2340 658 2540 734
use cut_M2M3_1x2 
transform 1 0 1912 0 1 596
box 1912 596 1988 796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1114
box 2340 1114 2540 1190
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1052
box 1912 1052 1988 1252
use cut_M1M3_2x1 
transform 1 0 2340 0 1 886
box 2340 886 2540 962
use cut_M2M3_1x2 
transform 1 0 1912 0 1 824
box 1912 824 1988 1024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 430
box 2340 430 2540 506
use cut_M2M3_1x2 
transform 1 0 1912 0 1 368
box 1912 368 1988 568
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1342
box 2340 1342 2540 1418
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1280
box 1912 1280 1988 1480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 658
box 2340 658 2540 734
use cut_M2M3_1x2 
transform 1 0 1912 0 1 596
box 1912 596 1988 796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1114
box 2340 1114 2540 1190
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1052
box 1912 1052 1988 1252
use cut_M1M3_2x1 
transform 1 0 2340 0 1 886
box 2340 886 2540 962
use cut_M2M3_1x2 
transform 1 0 1912 0 1 824
box 1912 824 1988 1024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 430
box 2340 430 2540 506
use cut_M2M3_1x2 
transform 1 0 1912 0 1 368
box 1912 368 1988 568
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1342
box 2340 1342 2540 1418
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1280
box 1912 1280 1988 1480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 658
box 2340 658 2540 734
use cut_M2M3_1x2 
transform 1 0 1912 0 1 596
box 1912 596 1988 796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1114
box 2340 1114 2540 1190
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1052
box 1912 1052 1988 1252
use cut_M1M3_2x1 
transform 1 0 2340 0 1 886
box 2340 886 2540 962
use cut_M2M3_1x2 
transform 1 0 1912 0 1 824
box 1912 824 1988 1024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 430
box 2340 430 2540 506
use cut_M2M3_1x2 
transform 1 0 1912 0 1 368
box 1912 368 1988 568
use cut_M1M3_2x1 
transform 1 0 2340 0 1 202
box 2340 202 2540 278
use cut_M2M3_1x2 
transform 1 0 1912 0 1 140
box 1912 140 1988 340
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1342
box 2340 1342 2540 1418
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1280
box 1912 1280 1988 1480
use cut_M1M3_2x1 
transform 1 0 2340 0 1 658
box 2340 658 2540 734
use cut_M2M3_1x2 
transform 1 0 1912 0 1 596
box 1912 596 1988 796
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1114
box 2340 1114 2540 1190
use cut_M2M3_1x2 
transform 1 0 1912 0 1 1052
box 1912 1052 1988 1252
use cut_M1M3_2x1 
transform 1 0 2340 0 1 886
box 2340 886 2540 962
use cut_M2M3_1x2 
transform 1 0 1912 0 1 824
box 1912 824 1988 1024
use cut_M1M3_2x1 
transform 1 0 2340 0 1 430
box 2340 430 2540 506
use cut_M2M3_1x2 
transform 1 0 1912 0 1 368
box 1912 368 1988 568
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6442
box 2340 6442 2540 6518
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6380
box 1912 6380 1988 6580
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7582
box 2340 7582 2540 7658
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7520
box 1912 7520 1988 7720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6898
box 2340 6898 2540 6974
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6836
box 1912 6836 1988 7036
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7354
box 2340 7354 2540 7430
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7292
box 1912 7292 1988 7492
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7126
box 2340 7126 2540 7202
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7064
box 1912 7064 1988 7264
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6670
box 2340 6670 2540 6746
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6608
box 1912 6608 1988 6808
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6442
box 2340 6442 2540 6518
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6380
box 1912 6380 1988 6580
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7582
box 2340 7582 2540 7658
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7520
box 1912 7520 1988 7720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6898
box 2340 6898 2540 6974
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6836
box 1912 6836 1988 7036
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7354
box 2340 7354 2540 7430
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7292
box 1912 7292 1988 7492
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7126
box 2340 7126 2540 7202
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7064
box 1912 7064 1988 7264
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6670
box 2340 6670 2540 6746
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6608
box 1912 6608 1988 6808
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6442
box 2340 6442 2540 6518
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6380
box 1912 6380 1988 6580
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7582
box 2340 7582 2540 7658
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7520
box 1912 7520 1988 7720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6898
box 2340 6898 2540 6974
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6836
box 1912 6836 1988 7036
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7354
box 2340 7354 2540 7430
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7292
box 1912 7292 1988 7492
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7126
box 2340 7126 2540 7202
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7064
box 1912 7064 1988 7264
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6670
box 2340 6670 2540 6746
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6608
box 1912 6608 1988 6808
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6442
box 2340 6442 2540 6518
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6380
box 1912 6380 1988 6580
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7582
box 2340 7582 2540 7658
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7520
box 1912 7520 1988 7720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6898
box 2340 6898 2540 6974
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6836
box 1912 6836 1988 7036
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7354
box 2340 7354 2540 7430
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7292
box 1912 7292 1988 7492
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7126
box 2340 7126 2540 7202
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7064
box 1912 7064 1988 7264
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6670
box 2340 6670 2540 6746
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6608
box 1912 6608 1988 6808
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6442
box 2340 6442 2540 6518
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6380
box 1912 6380 1988 6580
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7582
box 2340 7582 2540 7658
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7520
box 1912 7520 1988 7720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6898
box 2340 6898 2540 6974
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6836
box 1912 6836 1988 7036
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7354
box 2340 7354 2540 7430
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7292
box 1912 7292 1988 7492
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7126
box 2340 7126 2540 7202
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7064
box 1912 7064 1988 7264
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6670
box 2340 6670 2540 6746
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6608
box 1912 6608 1988 6808
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6442
box 2340 6442 2540 6518
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6380
box 1912 6380 1988 6580
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7582
box 2340 7582 2540 7658
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7520
box 1912 7520 1988 7720
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6898
box 2340 6898 2540 6974
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6836
box 1912 6836 1988 7036
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7354
box 2340 7354 2540 7430
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7292
box 1912 7292 1988 7492
use cut_M1M3_2x1 
transform 1 0 2340 0 1 7126
box 2340 7126 2540 7202
use cut_M2M3_1x2 
transform 1 0 1912 0 1 7064
box 1912 7064 1988 7264
use cut_M1M3_2x1 
transform 1 0 2340 0 1 6670
box 2340 6670 2540 6746
use cut_M2M3_1x2 
transform 1 0 1912 0 1 6608
box 1912 6608 1988 6808
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9562
box 2340 9562 2540 9638
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9500
box 1732 9500 1808 9700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10702
box 2340 10702 2540 10778
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10640
box 1732 10640 1808 10840
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10018
box 2340 10018 2540 10094
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9956
box 1732 9956 1808 10156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10474
box 2340 10474 2540 10550
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10412
box 1732 10412 1808 10612
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10246
box 2340 10246 2540 10322
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10184
box 1732 10184 1808 10384
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9790
box 2340 9790 2540 9866
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9728
box 1732 9728 1808 9928
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9562
box 2340 9562 2540 9638
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9500
box 1732 9500 1808 9700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10702
box 2340 10702 2540 10778
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10640
box 1732 10640 1808 10840
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10018
box 2340 10018 2540 10094
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9956
box 1732 9956 1808 10156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10474
box 2340 10474 2540 10550
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10412
box 1732 10412 1808 10612
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10246
box 2340 10246 2540 10322
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10184
box 1732 10184 1808 10384
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9790
box 2340 9790 2540 9866
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9728
box 1732 9728 1808 9928
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9562
box 2340 9562 2540 9638
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9500
box 1732 9500 1808 9700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10702
box 2340 10702 2540 10778
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10640
box 1732 10640 1808 10840
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10018
box 2340 10018 2540 10094
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9956
box 1732 9956 1808 10156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10474
box 2340 10474 2540 10550
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10412
box 1732 10412 1808 10612
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10246
box 2340 10246 2540 10322
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10184
box 1732 10184 1808 10384
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9790
box 2340 9790 2540 9866
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9728
box 1732 9728 1808 9928
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9562
box 2340 9562 2540 9638
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9500
box 1732 9500 1808 9700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10702
box 2340 10702 2540 10778
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10640
box 1732 10640 1808 10840
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10018
box 2340 10018 2540 10094
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9956
box 1732 9956 1808 10156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10474
box 2340 10474 2540 10550
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10412
box 1732 10412 1808 10612
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10246
box 2340 10246 2540 10322
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10184
box 1732 10184 1808 10384
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9790
box 2340 9790 2540 9866
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9728
box 1732 9728 1808 9928
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9562
box 2340 9562 2540 9638
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9500
box 1732 9500 1808 9700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10702
box 2340 10702 2540 10778
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10640
box 1732 10640 1808 10840
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10018
box 2340 10018 2540 10094
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9956
box 1732 9956 1808 10156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10474
box 2340 10474 2540 10550
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10412
box 1732 10412 1808 10612
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10246
box 2340 10246 2540 10322
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10184
box 1732 10184 1808 10384
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9790
box 2340 9790 2540 9866
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9728
box 1732 9728 1808 9928
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9562
box 2340 9562 2540 9638
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9500
box 1732 9500 1808 9700
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10702
box 2340 10702 2540 10778
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10640
box 1732 10640 1808 10840
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10018
box 2340 10018 2540 10094
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9956
box 1732 9956 1808 10156
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10474
box 2340 10474 2540 10550
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10412
box 1732 10412 1808 10612
use cut_M1M3_2x1 
transform 1 0 2340 0 1 10246
box 2340 10246 2540 10322
use cut_M2M3_1x2 
transform 1 0 1732 0 1 10184
box 1732 10184 1808 10384
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9790
box 2340 9790 2540 9866
use cut_M2M3_1x2 
transform 1 0 1732 0 1 9728
box 1732 9728 1808 9928
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1762
box 2340 1762 2540 1838
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1700
box 1552 1700 1628 1900
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2902
box 2340 2902 2540 2978
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2840
box 1552 2840 1628 3040
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2218
box 2340 2218 2540 2294
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2156
box 1552 2156 1628 2356
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2674
box 2340 2674 2540 2750
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2612
box 1552 2612 1628 2812
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2446
box 2340 2446 2540 2522
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2384
box 1552 2384 1628 2584
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1990
box 2340 1990 2540 2066
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1928
box 1552 1928 1628 2128
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1762
box 2340 1762 2540 1838
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1700
box 1552 1700 1628 1900
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2902
box 2340 2902 2540 2978
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2840
box 1552 2840 1628 3040
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2218
box 2340 2218 2540 2294
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2156
box 1552 2156 1628 2356
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2674
box 2340 2674 2540 2750
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2612
box 1552 2612 1628 2812
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2446
box 2340 2446 2540 2522
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2384
box 1552 2384 1628 2584
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1990
box 2340 1990 2540 2066
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1928
box 1552 1928 1628 2128
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1762
box 2340 1762 2540 1838
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1700
box 1552 1700 1628 1900
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2902
box 2340 2902 2540 2978
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2840
box 1552 2840 1628 3040
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2218
box 2340 2218 2540 2294
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2156
box 1552 2156 1628 2356
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2674
box 2340 2674 2540 2750
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2612
box 1552 2612 1628 2812
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2446
box 2340 2446 2540 2522
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2384
box 1552 2384 1628 2584
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1990
box 2340 1990 2540 2066
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1928
box 1552 1928 1628 2128
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1762
box 2340 1762 2540 1838
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1700
box 1552 1700 1628 1900
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2902
box 2340 2902 2540 2978
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2840
box 1552 2840 1628 3040
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2218
box 2340 2218 2540 2294
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2156
box 1552 2156 1628 2356
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2674
box 2340 2674 2540 2750
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2612
box 1552 2612 1628 2812
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2446
box 2340 2446 2540 2522
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2384
box 1552 2384 1628 2584
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1990
box 2340 1990 2540 2066
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1928
box 1552 1928 1628 2128
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1762
box 2340 1762 2540 1838
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1700
box 1552 1700 1628 1900
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2902
box 2340 2902 2540 2978
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2840
box 1552 2840 1628 3040
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2218
box 2340 2218 2540 2294
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2156
box 1552 2156 1628 2356
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2674
box 2340 2674 2540 2750
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2612
box 1552 2612 1628 2812
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2446
box 2340 2446 2540 2522
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2384
box 1552 2384 1628 2584
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1990
box 2340 1990 2540 2066
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1928
box 1552 1928 1628 2128
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1762
box 2340 1762 2540 1838
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1700
box 1552 1700 1628 1900
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2902
box 2340 2902 2540 2978
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2840
box 1552 2840 1628 3040
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2218
box 2340 2218 2540 2294
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2156
box 1552 2156 1628 2356
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2674
box 2340 2674 2540 2750
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2612
box 1552 2612 1628 2812
use cut_M1M3_2x1 
transform 1 0 2340 0 1 2446
box 2340 2446 2540 2522
use cut_M2M3_1x2 
transform 1 0 1552 0 1 2384
box 1552 2384 1628 2584
use cut_M1M3_2x1 
transform 1 0 2340 0 1 1990
box 2340 1990 2540 2066
use cut_M2M3_1x2 
transform 1 0 1552 0 1 1928
box 1552 1928 1628 2128
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3550
box 2340 3550 2540 3626
use cut_M2M3_1x2 
transform 1 0 1372 0 1 3488
box 1372 3488 1448 3688
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8230
box 2340 8230 2540 8306
use cut_M2M3_1x2 
transform 1 0 1192 0 1 8168
box 1192 8168 1268 8368
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8002
box 2340 8002 2540 8078
use cut_M2M3_1x2 
transform 1 0 1012 0 1 7940
box 1012 7940 1088 8140
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9142
box 2340 9142 2540 9218
use cut_M2M3_1x2 
transform 1 0 1012 0 1 9080
box 1012 9080 1088 9280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8458
box 2340 8458 2540 8534
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8396
box 1012 8396 1088 8596
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8914
box 2340 8914 2540 8990
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8852
box 1012 8852 1088 9052
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8002
box 2340 8002 2540 8078
use cut_M2M3_1x2 
transform 1 0 1012 0 1 7940
box 1012 7940 1088 8140
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9142
box 2340 9142 2540 9218
use cut_M2M3_1x2 
transform 1 0 1012 0 1 9080
box 1012 9080 1088 9280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8458
box 2340 8458 2540 8534
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8396
box 1012 8396 1088 8596
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8914
box 2340 8914 2540 8990
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8852
box 1012 8852 1088 9052
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8002
box 2340 8002 2540 8078
use cut_M2M3_1x2 
transform 1 0 1012 0 1 7940
box 1012 7940 1088 8140
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9142
box 2340 9142 2540 9218
use cut_M2M3_1x2 
transform 1 0 1012 0 1 9080
box 1012 9080 1088 9280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8458
box 2340 8458 2540 8534
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8396
box 1012 8396 1088 8596
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8914
box 2340 8914 2540 8990
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8852
box 1012 8852 1088 9052
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8002
box 2340 8002 2540 8078
use cut_M2M3_1x2 
transform 1 0 1012 0 1 7940
box 1012 7940 1088 8140
use cut_M1M3_2x1 
transform 1 0 2340 0 1 9142
box 2340 9142 2540 9218
use cut_M2M3_1x2 
transform 1 0 1012 0 1 9080
box 1012 9080 1088 9280
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8458
box 2340 8458 2540 8534
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8396
box 1012 8396 1088 8596
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8914
box 2340 8914 2540 8990
use cut_M2M3_1x2 
transform 1 0 1012 0 1 8852
box 1012 8852 1088 9052
use cut_M1M3_2x1 
transform 1 0 2340 0 1 8686
box 2340 8686 2540 8762
use cut_M2M3_1x2 
transform 1 0 832 0 1 8624
box 832 8624 908 8824
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4006
box 2340 4006 2540 4082
use cut_M2M3_1x2 
transform 1 0 652 0 1 3944
box 652 3944 728 4144
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4234
box 2340 4234 2540 4310
use cut_M2M3_1x2 
transform 1 0 472 0 1 4172
box 472 4172 548 4372
use cut_M1M3_2x1 
transform 1 0 2340 0 1 3778
box 2340 3778 2540 3854
use cut_M2M3_1x2 
transform 1 0 292 0 1 3716
box 292 3716 368 3916
use cut_M1M3_2x1 
transform 1 0 2340 0 1 4462
box 2340 4462 2540 4538
use cut_M2M3_1x2 
transform 1 0 112 0 1 4400
box 112 4400 188 4600
use cut_M1M2_1x2 
transform 1 0 2668 0 1 3268
box 2668 3268 2736 3452
use cut_M1M2_1x2 
transform 1 0 2668 0 1 3268
box 2668 3268 2736 3452
<< labels >>
flabel m1 s 2100 4820 2160 12480 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew
flabel m1 s 1920 140 1980 12480 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew
flabel m1 s 1740 9500 1800 12480 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew
flabel m1 s 1560 1700 1620 12480 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew
flabel m1 s 1380 3488 1440 12480 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew
flabel m1 s 1200 8168 1260 12480 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew
flabel m1 s 1020 7940 1080 12480 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew
flabel m1 s 840 8624 900 12480 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew
flabel m1 s 660 3944 720 12480 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew
flabel m1 s 480 4172 540 12480 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew
flabel m1 s 300 3716 360 12480 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew
flabel m1 s 120 4400 180 12480 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew
flabel m1 s 2668 0 11768 76 0 FreeSans 400 0 0 0 AVSS
port 14 nsew
flabel m3 s 2668 10920 2744 12540 0 FreeSans 400 0 0 0 CTOP
port 13 nsew
<< end >>
