magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 1920
<< locali >>
rect 360 770 514 830
rect 514 530 720 590
rect 514 530 574 830
rect 270 130 450 190
rect 270 450 450 510
rect 630 850 810 910
rect 2010 120 2190 200
rect -90 120 90 200
<< m3 >>
rect 1290 0 1474 1920
rect 630 0 814 1920
rect 1290 0 1474 1920
rect 630 0 814 1920
use NDX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2100 640
use IVX4_CV XA2
transform 1 0 0 0 1 640
box 0 640 2100 1920
<< labels >>
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 630 850 810 910 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel locali s 2010 120 2190 200 0 FreeSans 400 0 0 0 BULKP
port 4 nsew
flabel locali s -90 120 90 200 0 FreeSans 400 0 0 0 BULKN
port 5 nsew
flabel m3 s 1290 0 1474 1920 0 FreeSans 400 0 0 0 AVDD
port 6 nsew
flabel m3 s 630 0 814 1920 0 FreeSans 400 0 0 0 AVSS
port 7 nsew
<< end >>
