magic
tech sky130A
magscale 1 2
timestamp 1660233442
<< checkpaint >>
rect 0 0 68 184
<< locali >>
rect 0 0 68 184
<< viali >>
rect 6 12 62 68
rect 6 116 62 172
<< m1 >>
rect 0 0 68 184
<< labels >>
<< end >>
