magic
tech sky130A
magscale 1 2
timestamp 1658582973
<< checkpaint >>
rect 0 0 184 184
<< locali >>
rect 0 0 184 184
<< m1 >>
rect 0 0 184 184
<< viali >>
rect 12 12 172 172
<< labels >>
<< end >>
