magic
tech sky130A
magscale 1 2
timestamp 1660305041
<< checkpaint >>
rect 0 0 2520 1408
<< locali >>
rect 1626 234 1686 470
rect 1626 938 1686 1174
rect 1656 1290 1824 1350
rect 1824 498 2088 558
rect 1824 146 2088 206
rect 1824 146 1884 1350
rect 864 938 1032 998
rect 864 1290 1032 1350
rect 1032 938 1092 1350
rect 864 234 1032 294
rect 864 586 1032 646
rect 1032 234 1092 646
rect 432 146 600 206
rect 432 498 600 558
rect 600 146 660 558
rect 432 850 600 910
rect 432 1202 600 1262
rect 600 850 660 1262
rect 864 586 1032 646
rect 1032 586 1656 646
rect 1032 586 1092 646
rect 864 1290 1032 1350
rect 1032 1290 1656 1350
rect 1032 1290 1092 1350
rect 756 1290 972 1350
rect 324 850 540 910
rect 324 146 540 206
rect 756 234 972 294
<< m1 >>
rect 1656 586 1824 646
rect 1824 850 2088 910
rect 1824 1202 2088 1262
rect 1824 586 1884 1270
<< m3 >>
rect 1548 0 1748 1408
rect 756 0 956 1408
rect 1548 0 1748 1408
rect 756 0 956 1408
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xb1_00
transform 1 0 0 0 1 0
box 0 0 1260 352
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xb1_10
transform 1 0 0 0 1 352
box 0 352 1260 704
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xb2_00
transform 1 0 0 0 1 704
box 0 704 1260 1056
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xb2_10
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xc1a0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xc1b0
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xc2a0
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xc2b0
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use cut_M1M2_2x1 
transform 1 0 1548 0 1 586
box 1548 586 1732 654
use cut_M1M2_2x1 
transform 1 0 1980 0 1 850
box 1980 850 2164 918
use cut_M1M2_2x1 
transform 1 0 1980 0 1 1202
box 1980 1202 2164 1270
use cut_M1M4_2x1 
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use cut_M1M4_2x1 
transform 1 0 1548 0 1 762
box 1548 762 1748 838
use cut_M1M4_2x1 
transform 1 0 756 0 1 58
box 756 58 956 134
use cut_M1M4_2x1 
transform 1 0 756 0 1 410
box 756 410 956 486
use cut_M1M4_2x1 
transform 1 0 756 0 1 762
box 756 762 956 838
use cut_M1M4_2x1 
transform 1 0 756 0 1 1114
box 756 1114 956 1190
<< labels >>
flabel locali s 756 1290 972 1350 0 FreeSans 400 0 0 0 YN
port 3 nsew
flabel locali s 324 850 540 910 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 AN
port 2 nsew
flabel locali s 756 234 972 294 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel m3 s 1548 0 1748 1408 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 756 0 956 1408 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
