magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 184 184
<< m2 >>
rect 0 0 184 184
<< m3 >>
rect 0 0 184 184
<< v2 >>
rect 12 12 172 172
<< labels >>
<< end >>
