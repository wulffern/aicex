magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 1680 960
<< m1 >>
rect 120 -40 1640 40
rect 1560 40 1640 120
rect 120 120 1480 200
rect 1560 120 1640 200
rect 120 200 200 280
rect 1560 200 1640 280
rect 120 280 200 360
rect 280 280 1640 360
rect 120 360 200 440
rect 1560 360 1640 440
rect 120 440 1480 520
rect 1560 440 1640 520
rect 120 520 200 600
rect 1560 520 1640 600
rect 120 600 200 680
rect 280 600 1640 680
rect 120 680 200 760
rect 120 760 1640 840
<< m2 >>
rect 120 -40 1640 40
rect 1560 40 1640 120
rect 120 120 1480 200
rect 1560 120 1640 200
rect 120 200 200 280
rect 1560 200 1640 280
rect 120 280 200 360
rect 280 280 1640 360
rect 120 360 200 440
rect 1560 360 1640 440
rect 120 440 1480 520
rect 1560 440 1640 520
rect 120 520 200 600
rect 1560 520 1640 600
rect 120 600 200 680
rect 280 600 1640 680
rect 120 680 200 760
rect 120 760 1640 840
<< locali >>
rect 120 -40 1640 40
rect 1560 40 1640 120
rect 120 120 1480 200
rect 1560 120 1640 200
rect 120 200 200 280
rect 1560 200 1640 280
rect 120 280 200 360
rect 280 280 1640 360
rect 120 360 200 440
rect 1560 360 1640 440
rect 120 440 1480 520
rect 1560 440 1640 520
rect 120 520 200 600
rect 1560 520 1640 600
rect 120 600 200 680
rect 280 600 1640 680
rect 120 680 200 760
rect 120 760 1640 840
<< v1 >>
rect 1240 -32 1319 -24
rect 1240 -24 1319 -16
rect 1240 -16 1319 -8
rect 1240 -8 1319 0
rect 1240 0 1319 8
rect 1240 8 1319 16
rect 1240 16 1319 24
rect 1240 24 1319 32
rect 1320 -32 1399 -24
rect 1320 -24 1399 -16
rect 1320 -16 1399 -8
rect 1320 -8 1399 0
rect 1320 0 1399 8
rect 1320 8 1399 16
rect 1320 16 1399 24
rect 1320 24 1399 32
rect 1400 -32 1479 -24
rect 1400 -24 1479 -16
rect 1400 -16 1479 -8
rect 1400 -8 1479 0
rect 1400 0 1479 8
rect 1400 8 1479 16
rect 1400 16 1479 24
rect 1400 24 1479 32
rect 360 128 439 136
rect 360 136 439 144
rect 360 144 439 152
rect 360 152 439 160
rect 360 160 439 168
rect 360 168 439 176
rect 360 176 439 184
rect 360 184 439 192
rect 440 128 519 136
rect 440 136 519 144
rect 440 144 519 152
rect 440 152 519 160
rect 440 160 519 168
rect 440 168 519 176
rect 440 176 519 184
rect 440 184 519 192
rect 520 128 599 136
rect 520 136 599 144
rect 520 144 599 152
rect 520 152 599 160
rect 520 160 599 168
rect 520 168 599 176
rect 520 176 599 184
rect 520 184 599 192
rect 1240 288 1319 296
rect 1240 296 1319 304
rect 1240 304 1319 312
rect 1240 312 1319 320
rect 1240 320 1319 328
rect 1240 328 1319 336
rect 1240 336 1319 344
rect 1240 344 1319 352
rect 1320 288 1399 296
rect 1320 296 1399 304
rect 1320 304 1399 312
rect 1320 312 1399 320
rect 1320 320 1399 328
rect 1320 328 1399 336
rect 1320 336 1399 344
rect 1320 344 1399 352
rect 1400 288 1479 296
rect 1400 296 1479 304
rect 1400 304 1479 312
rect 1400 312 1479 320
rect 1400 320 1479 328
rect 1400 328 1479 336
rect 1400 336 1479 344
rect 1400 344 1479 352
rect 360 448 439 456
rect 360 456 439 464
rect 360 464 439 472
rect 360 472 439 480
rect 360 480 439 488
rect 360 488 439 496
rect 360 496 439 504
rect 360 504 439 512
rect 440 448 519 456
rect 440 456 519 464
rect 440 464 519 472
rect 440 472 519 480
rect 440 480 519 488
rect 440 488 519 496
rect 440 496 519 504
rect 440 504 519 512
rect 520 448 599 456
rect 520 456 599 464
rect 520 464 599 472
rect 520 472 599 480
rect 520 480 599 488
rect 520 488 599 496
rect 520 496 599 504
rect 520 504 599 512
rect 1240 608 1319 616
rect 1240 616 1319 624
rect 1240 624 1319 632
rect 1240 632 1319 640
rect 1240 640 1319 648
rect 1240 648 1319 656
rect 1240 656 1319 664
rect 1240 664 1319 672
rect 1320 608 1399 616
rect 1320 616 1399 624
rect 1320 624 1399 632
rect 1320 632 1399 640
rect 1320 640 1399 648
rect 1320 648 1399 656
rect 1320 656 1399 664
rect 1320 664 1399 672
rect 1400 608 1479 616
rect 1400 616 1479 624
rect 1400 624 1479 632
rect 1400 632 1479 640
rect 1400 640 1479 648
rect 1400 648 1479 656
rect 1400 656 1479 664
rect 1400 664 1479 672
rect 360 768 439 776
rect 360 776 439 784
rect 360 784 439 792
rect 360 792 439 800
rect 360 800 439 808
rect 360 808 439 816
rect 360 816 439 824
rect 360 824 439 832
rect 440 768 519 776
rect 440 776 519 784
rect 440 784 519 792
rect 440 792 519 800
rect 440 800 519 808
rect 440 808 519 816
rect 440 816 519 824
rect 440 824 519 832
rect 520 768 599 776
rect 520 776 599 784
rect 520 784 599 792
rect 520 792 599 800
rect 520 800 599 808
rect 520 808 599 816
rect 520 816 599 824
rect 520 824 599 832
<< v2 >>
rect 1240 -32 1319 -24
rect 1240 -24 1319 -16
rect 1240 -16 1319 -8
rect 1240 -8 1319 0
rect 1240 0 1319 8
rect 1240 8 1319 16
rect 1240 16 1319 24
rect 1240 24 1319 32
rect 1320 -32 1399 -24
rect 1320 -24 1399 -16
rect 1320 -16 1399 -8
rect 1320 -8 1399 0
rect 1320 0 1399 8
rect 1320 8 1399 16
rect 1320 16 1399 24
rect 1320 24 1399 32
rect 1400 -32 1479 -24
rect 1400 -24 1479 -16
rect 1400 -16 1479 -8
rect 1400 -8 1479 0
rect 1400 0 1479 8
rect 1400 8 1479 16
rect 1400 16 1479 24
rect 1400 24 1479 32
rect 360 128 439 136
rect 360 136 439 144
rect 360 144 439 152
rect 360 152 439 160
rect 360 160 439 168
rect 360 168 439 176
rect 360 176 439 184
rect 360 184 439 192
rect 440 128 519 136
rect 440 136 519 144
rect 440 144 519 152
rect 440 152 519 160
rect 440 160 519 168
rect 440 168 519 176
rect 440 176 519 184
rect 440 184 519 192
rect 520 128 599 136
rect 520 136 599 144
rect 520 144 599 152
rect 520 152 599 160
rect 520 160 599 168
rect 520 168 599 176
rect 520 176 599 184
rect 520 184 599 192
rect 1240 288 1319 296
rect 1240 296 1319 304
rect 1240 304 1319 312
rect 1240 312 1319 320
rect 1240 320 1319 328
rect 1240 328 1319 336
rect 1240 336 1319 344
rect 1240 344 1319 352
rect 1320 288 1399 296
rect 1320 296 1399 304
rect 1320 304 1399 312
rect 1320 312 1399 320
rect 1320 320 1399 328
rect 1320 328 1399 336
rect 1320 336 1399 344
rect 1320 344 1399 352
rect 1400 288 1479 296
rect 1400 296 1479 304
rect 1400 304 1479 312
rect 1400 312 1479 320
rect 1400 320 1479 328
rect 1400 328 1479 336
rect 1400 336 1479 344
rect 1400 344 1479 352
rect 360 448 439 456
rect 360 456 439 464
rect 360 464 439 472
rect 360 472 439 480
rect 360 480 439 488
rect 360 488 439 496
rect 360 496 439 504
rect 360 504 439 512
rect 440 448 519 456
rect 440 456 519 464
rect 440 464 519 472
rect 440 472 519 480
rect 440 480 519 488
rect 440 488 519 496
rect 440 496 519 504
rect 440 504 519 512
rect 520 448 599 456
rect 520 456 599 464
rect 520 464 599 472
rect 520 472 599 480
rect 520 480 599 488
rect 520 488 599 496
rect 520 496 599 504
rect 520 504 599 512
rect 1240 608 1319 616
rect 1240 616 1319 624
rect 1240 624 1319 632
rect 1240 632 1319 640
rect 1240 640 1319 648
rect 1240 648 1319 656
rect 1240 656 1319 664
rect 1240 664 1319 672
rect 1320 608 1399 616
rect 1320 616 1399 624
rect 1320 624 1399 632
rect 1320 632 1399 640
rect 1320 640 1399 648
rect 1320 648 1399 656
rect 1320 656 1399 664
rect 1320 664 1399 672
rect 1400 608 1479 616
rect 1400 616 1479 624
rect 1400 624 1479 632
rect 1400 632 1479 640
rect 1400 640 1479 648
rect 1400 648 1479 656
rect 1400 656 1479 664
rect 1400 664 1479 672
rect 360 768 439 776
rect 360 776 439 784
rect 360 784 439 792
rect 360 792 439 800
rect 360 800 439 808
rect 360 808 439 816
rect 360 816 439 824
rect 360 824 439 832
rect 440 768 519 776
rect 440 776 519 784
rect 440 784 519 792
rect 440 792 519 800
rect 440 800 519 808
rect 440 808 519 816
rect 440 816 519 824
rect 440 824 519 832
rect 520 768 599 776
rect 520 776 599 784
rect 520 784 599 792
rect 520 792 599 800
rect 520 800 599 808
rect 520 808 599 816
rect 520 816 599 824
rect 520 824 599 832
<< viali >>
rect 1240 -32 1319 -24
rect 1240 -24 1319 -16
rect 1240 -16 1319 -8
rect 1240 -8 1319 0
rect 1240 0 1319 8
rect 1240 8 1319 16
rect 1240 16 1319 24
rect 1240 24 1319 32
rect 1320 -32 1399 -24
rect 1320 -24 1399 -16
rect 1320 -16 1399 -8
rect 1320 -8 1399 0
rect 1320 0 1399 8
rect 1320 8 1399 16
rect 1320 16 1399 24
rect 1320 24 1399 32
rect 1400 -32 1479 -24
rect 1400 -24 1479 -16
rect 1400 -16 1479 -8
rect 1400 -8 1479 0
rect 1400 0 1479 8
rect 1400 8 1479 16
rect 1400 16 1479 24
rect 1400 24 1479 32
rect 360 128 439 136
rect 360 136 439 144
rect 360 144 439 152
rect 360 152 439 160
rect 360 160 439 168
rect 360 168 439 176
rect 360 176 439 184
rect 360 184 439 192
rect 440 128 519 136
rect 440 136 519 144
rect 440 144 519 152
rect 440 152 519 160
rect 440 160 519 168
rect 440 168 519 176
rect 440 176 519 184
rect 440 184 519 192
rect 520 128 599 136
rect 520 136 599 144
rect 520 144 599 152
rect 520 152 599 160
rect 520 160 599 168
rect 520 168 599 176
rect 520 176 599 184
rect 520 184 599 192
rect 1240 288 1319 296
rect 1240 296 1319 304
rect 1240 304 1319 312
rect 1240 312 1319 320
rect 1240 320 1319 328
rect 1240 328 1319 336
rect 1240 336 1319 344
rect 1240 344 1319 352
rect 1320 288 1399 296
rect 1320 296 1399 304
rect 1320 304 1399 312
rect 1320 312 1399 320
rect 1320 320 1399 328
rect 1320 328 1399 336
rect 1320 336 1399 344
rect 1320 344 1399 352
rect 1400 288 1479 296
rect 1400 296 1479 304
rect 1400 304 1479 312
rect 1400 312 1479 320
rect 1400 320 1479 328
rect 1400 328 1479 336
rect 1400 336 1479 344
rect 1400 344 1479 352
rect 360 448 439 456
rect 360 456 439 464
rect 360 464 439 472
rect 360 472 439 480
rect 360 480 439 488
rect 360 488 439 496
rect 360 496 439 504
rect 360 504 439 512
rect 440 448 519 456
rect 440 456 519 464
rect 440 464 519 472
rect 440 472 519 480
rect 440 480 519 488
rect 440 488 519 496
rect 440 496 519 504
rect 440 504 519 512
rect 520 448 599 456
rect 520 456 599 464
rect 520 464 599 472
rect 520 472 599 480
rect 520 480 599 488
rect 520 488 599 496
rect 520 496 599 504
rect 520 504 599 512
rect 1240 608 1319 616
rect 1240 616 1319 624
rect 1240 624 1319 632
rect 1240 632 1319 640
rect 1240 640 1319 648
rect 1240 648 1319 656
rect 1240 656 1319 664
rect 1240 664 1319 672
rect 1320 608 1399 616
rect 1320 616 1399 624
rect 1320 624 1399 632
rect 1320 632 1399 640
rect 1320 640 1399 648
rect 1320 648 1399 656
rect 1320 656 1399 664
rect 1320 664 1399 672
rect 1400 608 1479 616
rect 1400 616 1479 624
rect 1400 624 1479 632
rect 1400 632 1479 640
rect 1400 640 1479 648
rect 1400 648 1479 656
rect 1400 656 1479 664
rect 1400 664 1479 672
rect 360 768 439 776
rect 360 776 439 784
rect 360 784 439 792
rect 360 792 439 800
rect 360 800 439 808
rect 360 808 439 816
rect 360 816 439 824
rect 360 824 439 832
rect 440 768 519 776
rect 440 776 519 784
rect 440 784 519 792
rect 440 792 519 800
rect 440 800 519 808
rect 440 808 519 816
rect 440 816 519 824
rect 440 824 519 832
rect 520 768 599 776
rect 520 776 599 784
rect 520 784 599 792
rect 520 792 599 800
rect 520 800 599 808
rect 520 808 599 816
rect 520 816 599 824
rect 520 824 599 832
<< m3 >>
rect 120 -40 1640 40
rect 1560 40 1640 120
rect 120 120 1240 200
rect 1320 120 1480 200
rect 1560 120 1640 200
rect 120 200 200 280
rect 1560 200 1640 280
rect 120 280 200 360
rect 280 280 360 360
rect 440 280 1640 360
rect 120 360 200 440
rect 1560 360 1640 440
rect 120 440 1480 520
rect 1560 440 1640 520
rect 120 520 200 600
rect 1560 520 1640 600
rect 120 600 200 680
rect 280 600 1640 680
rect 120 680 200 760
rect 120 760 1640 840
<< rm3 >>
rect 1240 120 1320 200
rect 360 280 440 360
<< labels >>
flabel m3 s 120 -40 1640 40 0 FreeSans 400 0 0 0 B
port 1 nsew
flabel m3 s 120 760 1640 840 0 FreeSans 400 0 0 0 A
port 2 nsew
<< end >>
