magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 1600
<< locali >>
rect 720 210 874 270
rect 720 370 874 430
rect 720 690 874 750
rect 720 1010 874 1070
rect 874 210 934 1070
rect 1166 210 1380 270
rect 1166 370 1380 430
rect 1166 850 1380 910
rect 1166 1170 1380 1230
rect 1166 210 1226 1230
rect 330 130 390 510
rect 1740 770 1894 830
rect 1380 530 1894 590
rect 1740 1090 1894 1150
rect 1740 1410 1894 1470
rect 1894 530 1954 1470
rect 146 770 360 830
rect 146 530 720 590
rect 146 1090 360 1150
rect 146 1410 360 1470
rect 146 530 206 1470
rect 506 850 720 910
rect 506 1170 720 1230
rect 506 850 566 1230
rect 720 1490 874 1550
rect 874 1490 1380 1550
rect 874 1490 934 1550
rect 720 1170 874 1230
rect 874 1330 1380 1390
rect 874 1170 934 1390
rect 1380 690 1534 750
rect 1380 1010 1534 1070
rect 1534 690 1594 1070
rect 270 130 450 190
rect 630 1490 810 1550
<< m1 >>
rect 720 1330 874 1390
rect 874 1010 1380 1070
rect 874 1010 934 1398
rect 720 530 874 590
rect 874 530 1380 590
rect 874 530 934 598
<< poly >>
rect 270 142 1830 178
rect 270 462 1830 498
<< m3 >>
rect 1290 0 1474 1600
rect 630 0 814 1600
rect 1290 0 1474 1600
rect 630 0 814 1600
use NCHDL XA2
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL XA3
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL XA4a
transform 1 0 0 0 1 640
box 0 640 1050 960
use NCHDL XA4b
transform 1 0 0 0 1 960
box 0 960 1050 1280
use NCHDL XA5
transform 1 0 0 0 1 1280
box 0 1280 1050 1600
use PCHDL XB0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL XB1
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL XB3a
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use PCHDL XB3b
transform 1 0 1050 0 1 960
box 1050 960 2100 1280
use PCHDL XB4
transform 1 0 1050 0 1 1280
box 1050 1280 2100 1600
use cut_M1M2_2x1 
transform 1 0 630 0 1 1330
box 630 1330 814 1398
use cut_M1M2_2x1 
transform 1 0 1290 0 1 1010
box 1290 1010 1474 1078
use cut_M1M2_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M2_2x1 
transform 1 0 1290 0 1 530
box 1290 530 1474 598
use cut_M1M4_2x1 
transform 1 0 1290 0 1 50
box 1290 50 1474 118
use cut_M1M4_2x1 
transform 1 0 1290 0 1 1330
box 1290 1330 1474 1398
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 1330
box 630 1330 814 1398
<< labels >>
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 630 1490 810 1550 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel m3 s 1290 0 1474 1600 0 FreeSans 400 0 0 0 AVDD
port 3 nsew
flabel m3 s 630 0 814 1600 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
<< end >>
