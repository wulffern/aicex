magic
tech sky130A
magscale 1 2
timestamp 1658600916
<< checkpaint >>
rect -2284 0 26372 40022
<< m3 >>
rect 9100 18520 26178 18596
rect 9100 18908 26178 18984
rect 24104 19288 24180 26792
rect 24384 19288 24460 34536
rect 3944 19372 4020 30304
rect 4824 19566 4900 30304
rect 8984 19760 9060 30304
rect -216 19954 -140 30304
rect -216 19954 -140 30304
rect 13432 20148 13508 30330
rect 13432 20148 13508 30330
rect 18472 20342 18548 30330
rect 18472 20342 18548 30330
rect 10579 20536 10655 30330
rect 10579 20536 10655 30330
rect 15619 20730 15695 30330
rect 15619 20730 15695 30330
rect 499 20924 575 30330
rect 5539 21118 5615 30330
rect 5539 21118 5615 30330
rect 3352 21312 3428 30330
rect 3352 21312 3428 30330
rect 8392 21506 8468 30330
rect 8392 21506 8468 30330
rect 659 21700 735 31738
rect 8232 21894 8308 31738
rect 5699 22088 5775 31738
rect 3192 22282 3268 31738
rect 10914 22476 10990 33146
rect 13098 22670 13174 33146
rect 15954 22864 16030 33146
rect 8058 23058 8134 33146
rect 3018 23252 3094 33146
rect 834 23446 910 33146
rect 18138 23640 18214 33146
rect 5874 23834 5950 33146
rect 11072 50 11272 126
rect 12816 50 13016 126
rect 20659 30330 20735 30530
rect 1568 29344 1768 29544
rect 8856 0 9056 5280
rect 9648 0 9848 5280
<< m2 >>
rect 14872 18014 14948 18596
rect 9100 18014 9176 18984
rect 3944 19296 14020 19372
rect 4824 19490 13660 19566
rect 8984 19684 13300 19760
rect -216 19878 14380 19954
rect 11304 20072 13508 20148
rect 11664 20266 18548 20342
rect 10579 20460 11200 20536
rect 11484 20654 15695 20730
rect 499 20848 9760 20924
rect 5539 21042 10480 21118
rect 3352 21236 10120 21312
rect 8392 21430 10840 21506
rect 659 21624 9940 21700
rect 8232 21818 11020 21894
rect 5699 22012 10660 22088
rect 3192 22206 10300 22282
rect 10914 22400 12940 22476
rect 12684 22594 13174 22670
rect 12504 22788 16030 22864
rect 8058 22982 13120 23058
rect 3018 23176 13840 23252
rect 834 23370 14200 23446
rect 12324 23564 18214 23640
rect 5874 23758 13480 23834
rect -216 25024 -16 25100
<< m4 >>
rect 24104 18908 24180 19288
rect 24384 18520 24460 19288
<< m1 >>
rect 13944 17954 14020 19296
rect 13584 17954 13660 19490
rect 13224 17954 13300 19684
rect 14304 17954 14380 19878
rect 11304 17954 11380 20072
rect 11664 17954 11740 20266
rect 11124 17954 11200 20460
rect 11484 17954 11560 20654
rect 9684 17954 9760 20848
rect 10404 17954 10480 21042
rect 10044 17954 10120 21236
rect 10764 17954 10840 21430
rect 9864 17954 9940 21624
rect 10944 17954 11020 21818
rect 10584 17954 10660 22012
rect 10224 17954 10300 22206
rect 12864 17954 12940 22400
rect 12684 17954 12760 22594
rect 12504 17954 12580 22788
rect 13044 17954 13120 22982
rect 13764 17954 13840 23176
rect 14124 17954 14200 23370
rect 12324 17954 12400 23564
rect 13404 17954 13480 23758
<< locali >>
rect 11072 2698 11288 2758
rect 11072 1290 11288 1350
rect 20360 36384 20576 36444
rect -232 34888 -16 34948
rect 10064 498 10280 558
use SARBSSW_CV XB1
transform -1 0 12044 0 1 0
box 12044 0 26372 5280
use SARBSSW_CV XB2
transform 1 0 12044 0 1 0
box 12044 0 26372 5280
use CDAC8_CV XDAC1
transform -1 0 11844 0 1 5474
box 11844 5474 23576 18014
use CDAC8_CV XDAC2
transform 1 0 12204 0 1 5474
box 12204 5474 23936 18014
use SARDIGEX4_CV XA0
transform 1 0 -556 0 1 24534
box -556 24534 1964 38966
use SARDIGEX4_CV XA1
transform -1 0 4484 0 1 24534
box 4484 24534 7004 38966
use SARDIGEX4_CV XA2
transform 1 0 4484 0 1 24534
box 4484 24534 7004 38966
use SARDIGEX4_CV XA3
transform -1 0 9524 0 1 24534
box 9524 24534 12044 38966
use SARDIGEX4_CV XA4
transform 1 0 9524 0 1 24534
box 9524 24534 12044 38966
use SARDIGEX4_CV XA5
transform -1 0 14564 0 1 24534
box 14564 24534 17084 38966
use SARDIGEX4_CV XA6
transform 1 0 14564 0 1 24534
box 14564 24534 17084 38966
use SARDIGEX4_CV XA7
transform -1 0 19604 0 1 24534
box 19604 24534 22124 38966
use SARDIGEX4_CV XA8
transform 1 0 19604 0 1 24534
box 19604 24534 22124 38966
use SARCMPX1_CV XA20
transform -1 0 24644 0 1 24534
box 24644 24534 27164 40022
use cut_M3M4_1x2 
transform 1 0 14872 0 1 18014
box 14872 18014 14948 18214
use cut_M3M4_2x1 
transform 1 0 14872 0 1 18520
box 14872 18520 15072 18596
use cut_M3M4_1x2 
transform 1 0 9100 0 1 18014
box 9100 18014 9176 18214
use cut_M3M4_2x1 
transform 1 0 9100 0 1 18908
box 9100 18908 9300 18984
use cut_M2M4_2x1 
transform 1 0 24104 0 1 26792
box 24104 26792 24304 26868
use cut_M4M5_2x1 
transform 1 0 24104 0 1 18908
box 24104 18908 24304 18984
use cut_M4M5_1x2 
transform 1 0 24104 0 1 19288
box 24104 19288 24180 19488
use cut_M3M4_2x1 
transform 1 0 24260 0 1 34536
box 24260 34536 24460 34612
use cut_M2M3_2x1 
transform 1 0 24104 0 1 34536
box 24104 34536 24304 34612
use cut_M4M5_2x1 
transform 1 0 24384 0 1 18520
box 24384 18520 24584 18596
use cut_M4M5_1x2 
transform 1 0 24384 0 1 19288
box 24384 19288 24460 19488
use cut_M3M4_1x2 
transform 1 0 3944 0 1 19234
box 3944 19234 4020 19434
use cut_M2M3_1x2 
transform 1 0 13936 0 1 19234
box 13936 19234 14012 19434
use cut_M3M4_1x2 
transform 1 0 4824 0 1 19428
box 4824 19428 4900 19628
use cut_M2M3_1x2 
transform 1 0 13576 0 1 19428
box 13576 19428 13652 19628
use cut_M3M4_1x2 
transform 1 0 8984 0 1 19622
box 8984 19622 9060 19822
use cut_M2M3_1x2 
transform 1 0 13216 0 1 19622
box 13216 19622 13292 19822
use cut_M3M4_1x2 
transform 1 0 -216 0 1 19816
box -216 19816 -140 20016
use cut_M2M3_1x2 
transform 1 0 14296 0 1 19816
box 14296 19816 14372 20016
use cut_M3M4_1x2 
transform 1 0 13432 0 1 20010
box 13432 20010 13508 20210
use cut_M2M3_1x2 
transform 1 0 11296 0 1 20010
box 11296 20010 11372 20210
use cut_M3M4_1x2 
transform 1 0 18472 0 1 20204
box 18472 20204 18548 20404
use cut_M2M3_1x2 
transform 1 0 11656 0 1 20204
box 11656 20204 11732 20404
use cut_M3M4_1x2 
transform 1 0 10579 0 1 20398
box 10579 20398 10655 20598
use cut_M2M3_1x2 
transform 1 0 11116 0 1 20398
box 11116 20398 11192 20598
use cut_M3M4_1x2 
transform 1 0 15619 0 1 20592
box 15619 20592 15695 20792
use cut_M2M3_1x2 
transform 1 0 11476 0 1 20592
box 11476 20592 11552 20792
use cut_M3M4_1x2 
transform 1 0 499 0 1 20786
box 499 20786 575 20986
use cut_M2M3_1x2 
transform 1 0 9676 0 1 20786
box 9676 20786 9752 20986
use cut_M3M4_1x2 
transform 1 0 5539 0 1 20980
box 5539 20980 5615 21180
use cut_M2M3_1x2 
transform 1 0 10396 0 1 20980
box 10396 20980 10472 21180
use cut_M3M4_1x2 
transform 1 0 3352 0 1 21174
box 3352 21174 3428 21374
use cut_M2M3_1x2 
transform 1 0 10036 0 1 21174
box 10036 21174 10112 21374
use cut_M3M4_1x2 
transform 1 0 8392 0 1 21368
box 8392 21368 8468 21568
use cut_M2M3_1x2 
transform 1 0 10756 0 1 21368
box 10756 21368 10832 21568
use cut_M3M4_1x2 
transform 1 0 659 0 1 21562
box 659 21562 735 21762
use cut_M2M3_1x2 
transform 1 0 9856 0 1 21562
box 9856 21562 9932 21762
use cut_M3M4_1x2 
transform 1 0 8232 0 1 21756
box 8232 21756 8308 21956
use cut_M2M3_1x2 
transform 1 0 10936 0 1 21756
box 10936 21756 11012 21956
use cut_M3M4_1x2 
transform 1 0 5699 0 1 21950
box 5699 21950 5775 22150
use cut_M2M3_1x2 
transform 1 0 10576 0 1 21950
box 10576 21950 10652 22150
use cut_M3M4_1x2 
transform 1 0 3192 0 1 22144
box 3192 22144 3268 22344
use cut_M2M3_1x2 
transform 1 0 10216 0 1 22144
box 10216 22144 10292 22344
use cut_M3M4_1x2 
transform 1 0 10914 0 1 22338
box 10914 22338 10990 22538
use cut_M2M3_1x2 
transform 1 0 12856 0 1 22338
box 12856 22338 12932 22538
use cut_M3M4_1x2 
transform 1 0 13098 0 1 22532
box 13098 22532 13174 22732
use cut_M2M3_1x2 
transform 1 0 12676 0 1 22532
box 12676 22532 12752 22732
use cut_M3M4_1x2 
transform 1 0 15954 0 1 22726
box 15954 22726 16030 22926
use cut_M2M3_1x2 
transform 1 0 12496 0 1 22726
box 12496 22726 12572 22926
use cut_M3M4_1x2 
transform 1 0 8058 0 1 22920
box 8058 22920 8134 23120
use cut_M2M3_1x2 
transform 1 0 13036 0 1 22920
box 13036 22920 13112 23120
use cut_M3M4_1x2 
transform 1 0 3018 0 1 23114
box 3018 23114 3094 23314
use cut_M2M3_1x2 
transform 1 0 13756 0 1 23114
box 13756 23114 13832 23314
use cut_M3M4_1x2 
transform 1 0 834 0 1 23308
box 834 23308 910 23508
use cut_M2M3_1x2 
transform 1 0 14116 0 1 23308
box 14116 23308 14192 23508
use cut_M3M4_1x2 
transform 1 0 18138 0 1 23502
box 18138 23502 18214 23702
use cut_M2M3_1x2 
transform 1 0 12316 0 1 23502
box 12316 23502 12392 23702
use cut_M3M4_1x2 
transform 1 0 5874 0 1 23696
box 5874 23696 5950 23896
use cut_M2M3_1x2 
transform 1 0 13396 0 1 23696
box 13396 23696 13472 23896
<< labels >>
flabel m3 s -216 19954 -140 30304 0 FreeSans 400 0 0 0 D<8>
port 6 nsew
flabel m3 s 13432 20148 13508 30330 0 FreeSans 400 0 0 0 D<3>
port 11 nsew
flabel m3 s 18472 20342 18548 30330 0 FreeSans 400 0 0 0 D<1>
port 13 nsew
flabel m3 s 10579 20536 10655 30330 0 FreeSans 400 0 0 0 D<4>
port 10 nsew
flabel m3 s 15619 20730 15695 30330 0 FreeSans 400 0 0 0 D<2>
port 12 nsew
flabel m3 s 5539 21118 5615 30330 0 FreeSans 400 0 0 0 D<6>
port 8 nsew
flabel m3 s 3352 21312 3428 30330 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8392 21506 8468 30330 0 FreeSans 400 0 0 0 D<5>
port 9 nsew
flabel m3 s 11072 50 11272 126 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew
flabel m3 s 12816 50 13016 126 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew
flabel locali s 11072 2698 11288 2758 0 FreeSans 400 0 0 0 SARN
port 3 nsew
flabel locali s 11072 1290 11288 1350 0 FreeSans 400 0 0 0 SARP
port 4 nsew
flabel locali s 20360 36384 20576 36444 0 FreeSans 400 0 0 0 DONE
port 5 nsew
flabel m3 s 20659 30330 20735 30530 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
flabel m2 s -216 25024 -16 25100 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s -232 34888 -16 34948 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 10064 498 10280 558 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel m3 s 1568 29344 1768 29544 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel m3 s 8856 0 9056 5280 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel m3 s 9648 0 9848 5280 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
<< end >>
