** sch_path: /Users/wulff/pro/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_ROSC.sch
**.subckt SUN_PLL_ROSC PWRUP_1V8 VDD_ROSC AVSS VDD_1V8 CK
*.iopin PWRUP_1V8
*.iopin VDD_ROSC
*.iopin AVSS
*.iopin VDD_1V8
*.iopin CK
x1[7] AVSS VDD_ROSC NI N[7] SUNTR_IVX1_CV
x1[6] AVSS VDD_ROSC N[7] N[6] SUNTR_IVX1_CV
x1[5] AVSS VDD_ROSC N[6] N[5] SUNTR_IVX1_CV
x1[4] AVSS VDD_ROSC N[5] N[4] SUNTR_IVX1_CV
x1[3] AVSS VDD_ROSC N[4] N[3] SUNTR_IVX1_CV
x1[2] AVSS VDD_ROSC N[3] N[2] SUNTR_IVX1_CV
x1[1] AVSS VDD_ROSC N[2] N[1] SUNTR_IVX1_CV
x1[0] AVSS VDD_ROSC N[1] N[0] SUNTR_IVX1_CV
x1 AVSS VDD_ROSC N[0] PWRUP_1V8 NI SUNTR_NDX1_CV
x2 net1 CKUP VDD_1V8 VDD_1V8 SUNTR_PCHDL
x3 CKUP net1 VDD_1V8 VDD_1V8 SUNTR_PCHDL
x4 N[1] CKUP AVSS AVSS SUNTR_NCHDLA
x5 N[0] net1 AVSS AVSS SUNTR_NCHDLA
x6 AVSS VDD_1V8 CKUP CK SUNTR_IVX1_CV
**.ends

* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_IVX1_CV.sym # of pins=4
** sym_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV.sym
** sch_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV.sch
.subckt SUNTR_IVX1_CV  AVSS AVDD A Y
*.ipin A
*.opin Y
*.ipin AVDD
*.ipin AVSS
XMN0 A Y AVSS AVSS SUNTR_NCHDL
XMP0 A Y AVDD AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NDX1_CV.sym # of pins=5
** sym_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NDX1_CV.sym
** sch_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NDX1_CV.sch
.subckt SUNTR_NDX1_CV  AVSS AVDD B A Y
*.iopin A
*.iopin B
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 A N1 AVSS AVSS SUNTR_NCHDL
XMN1 B Y AVSS N1 SUNTR_NCHDL
XMP0 A Y AVDD AVDD SUNTR_PCHDL
XMP1 B AVDD AVDD Y SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_PCHDL.sym # of pins=4
** sym_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL.sym
** sch_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL.sch
.subckt SUNTR_PCHDL  G D B S
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.18 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHDLA.sym # of pins=4
** sym_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA.sym
** sch_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA.sch
.subckt SUNTR_NCHDLA  G D B S
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0 G D B S SUNTR_NCHDL
XM1 G S B D SUNTR_NCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHDL.sym # of pins=4
** sym_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL.sym
** sch_path: /Users/wulff/pro/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL.sch
.subckt SUNTR_NCHDL  G D B S
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.18 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
