magic
tech sky130A
magscale 1 2
timestamp 1658600916
<< checkpaint >>
rect 0 30 9504 1590
<< m3 >>
rect 328 0 404 1620
rect 328 0 404 1620
rect 468 140 544 1480
rect 608 0 684 1620
rect 748 140 824 1480
rect 888 0 964 1620
rect 1028 140 1104 1480
rect 1168 0 1244 1620
rect 1308 140 1384 1480
rect 1448 0 1524 1620
rect 1588 140 1664 1480
rect 1728 0 1804 1620
rect 1868 140 1944 1480
rect 2008 0 2084 1620
rect 2148 140 2224 1480
rect 2288 0 2364 1620
rect 2428 140 2504 1480
rect 2568 0 2644 1620
rect 2708 140 2784 1480
rect 2848 0 2924 1620
rect 2988 140 3064 1480
rect 3128 0 3204 1620
rect 3268 140 3344 1480
rect 3408 0 3484 1620
rect 3548 140 3624 1480
rect 3688 0 3764 1620
rect 3828 140 3904 1480
rect 3968 0 4044 1620
rect 4108 140 4184 1480
rect 4248 0 4324 1620
rect 4388 140 4464 1480
rect 4528 0 4604 1620
rect 4668 140 4744 1480
rect 4808 0 4884 1620
rect 4948 140 5024 1480
rect 5088 0 5164 1620
rect 5228 140 5304 1480
rect 5368 0 5444 1620
rect 5508 140 5584 1480
rect 5648 0 5724 1620
rect 5788 140 5864 1480
rect 5928 0 6004 1620
rect 6068 140 6144 1480
rect 6208 0 6284 1620
rect 6348 140 6424 1480
rect 6488 0 6564 1620
rect 6628 140 6704 1480
rect 6768 0 6844 1620
rect 6908 140 6984 1480
rect 7048 0 7124 1620
rect 7188 140 7264 1480
rect 7328 0 7404 1620
rect 7468 140 7544 1480
rect 7608 0 7684 1620
rect 7748 140 7824 1480
rect 7888 0 7964 1620
rect 8028 140 8104 1480
rect 8168 0 8244 1620
rect 8308 140 8384 1480
rect 8448 0 8524 1620
rect 8588 140 8664 1480
rect 8728 0 8804 1620
rect 8868 140 8944 1480
rect 9008 0 9084 1620
rect 9148 140 9224 1480
rect 9428 0 9504 1620
rect 9288 0 9364 1620
rect 328 0 9288 76
rect 328 1544 9288 1620
<< m1 >>
rect 328 0 9428 76
rect 2428 400 2504 1620
rect 7188 0 7264 1220
rect 2708 0 2784 536
rect 2708 856 2784 1620
rect 6908 0 6984 536
rect 6908 856 6984 1620
rect 2148 0 2224 992
rect 2148 1312 2224 1620
rect 2988 0 3064 992
rect 2988 1312 3064 1620
rect 6628 0 6704 992
rect 6628 1312 6704 1620
rect 7468 0 7544 992
rect 7468 1312 7544 1620
rect 1588 0 1664 764
rect 1588 1084 1664 1620
rect 1868 0 1944 764
rect 1868 1084 1944 1620
rect 3268 0 3344 764
rect 3268 1084 3344 1620
rect 3548 0 3624 764
rect 3548 1084 3624 1620
rect 6068 0 6144 764
rect 6068 1084 6144 1620
rect 6348 0 6424 764
rect 6348 1084 6424 1620
rect 7748 0 7824 764
rect 7748 1084 7824 1620
rect 8028 0 8104 764
rect 8028 1084 8104 1620
rect 468 0 544 308
rect 468 628 544 1620
rect 748 0 824 308
rect 748 628 824 1620
rect 1028 0 1104 308
rect 1028 628 1104 1620
rect 1308 0 1384 308
rect 1308 628 1384 1620
rect 3828 0 3904 308
rect 3828 628 3904 1620
rect 4108 0 4184 308
rect 4108 628 4184 1620
rect 4388 0 4464 308
rect 4388 628 4464 1620
rect 4668 0 4744 308
rect 4668 628 4744 1620
rect 4948 0 5024 308
rect 4948 628 5024 1620
rect 5228 0 5304 308
rect 5228 628 5304 1620
rect 5508 0 5584 308
rect 5508 628 5584 1620
rect 5788 0 5864 308
rect 5788 628 5864 1620
rect 8308 0 8384 308
rect 8308 628 8384 1620
rect 8588 0 8664 308
rect 8588 628 8664 1620
rect 8868 0 8944 308
rect 8868 628 8944 1620
rect 9148 0 9224 308
rect 9148 628 9224 1620
rect 328 0 404 1544
rect 608 0 684 1544
rect 888 0 964 1544
rect 1168 0 1244 1544
rect 1448 0 1524 1544
rect 1728 0 1804 1544
rect 2008 0 2084 1544
rect 2288 0 2364 1544
rect 2568 0 2644 1544
rect 2848 0 2924 1544
rect 3128 0 3204 1544
rect 3408 0 3484 1544
rect 3688 0 3764 1544
rect 3968 0 4044 1544
rect 4248 0 4324 1544
rect 4528 0 4604 1544
rect 4808 0 4884 1544
rect 5088 0 5164 1544
rect 5368 0 5444 1544
rect 5648 0 5724 1544
rect 5928 0 6004 1544
rect 6208 0 6284 1544
rect 6488 0 6564 1544
rect 6768 0 6844 1544
rect 7048 0 7124 1544
rect 7328 0 7404 1544
rect 7608 0 7684 1544
rect 7888 0 7964 1544
rect 8168 0 8244 1544
rect 8448 0 8524 1544
rect 8728 0 8804 1544
rect 9008 0 9084 1544
rect 9428 0 9504 1620
rect 9288 0 9364 1620
rect 328 0 9428 76
rect 328 1544 9428 1620
<< locali >>
rect 0 202 200 278
rect 0 1342 200 1418
rect 0 658 200 734
rect 0 1114 200 1190
rect 0 886 200 962
rect 0 430 200 506
rect 320 430 9288 506
rect 320 202 9288 278
rect 320 1342 9288 1418
rect 320 658 9288 734
rect 320 1114 9288 1190
rect 320 886 9288 962
<< m4 >>
rect 188 0 264 1620
rect 468 0 544 1620
rect 748 0 824 1620
rect 1028 0 1104 1620
rect 1308 0 1384 1620
rect 1588 0 1664 1620
rect 1868 0 1944 1620
rect 2148 0 2224 1620
rect 2428 0 2504 1620
rect 2708 0 2784 1620
rect 2988 0 3064 1620
rect 3268 0 3344 1620
rect 3548 0 3624 1620
rect 3828 0 3904 1620
rect 4108 0 4184 1620
rect 4388 0 4464 1620
rect 4668 0 4744 1620
rect 4948 0 5024 1620
rect 5228 0 5304 1620
rect 5508 0 5584 1620
rect 5788 0 5864 1620
rect 6068 0 6144 1620
rect 6348 0 6424 1620
rect 6628 0 6704 1620
rect 6908 0 6984 1620
rect 7188 0 7264 1620
rect 7468 0 7544 1620
rect 7748 0 7824 1620
rect 8028 0 8104 1620
rect 8308 0 8384 1620
rect 8588 0 8664 1620
rect 8868 0 8944 1620
rect 9148 0 9224 1620
rect 9428 0 9504 1620
rect 188 0 9428 76
rect 188 1544 9428 1620
<< m2 >>
rect 468 140 544 1480
rect 748 140 824 1480
rect 1028 140 1104 1480
rect 1308 140 1384 1480
rect 1588 140 1664 1480
rect 1868 140 1944 1480
rect 2148 140 2224 1480
rect 2428 140 2504 1480
rect 2708 140 2784 1480
rect 2988 140 3064 1480
rect 3268 140 3344 1480
rect 3548 140 3624 1480
rect 3828 140 3904 1480
rect 4108 140 4184 1480
rect 4388 140 4464 1480
rect 4668 140 4744 1480
rect 4948 140 5024 1480
rect 5228 140 5304 1480
rect 5508 140 5584 1480
rect 5788 140 5864 1480
rect 6068 140 6144 1480
rect 6348 140 6424 1480
rect 6628 140 6704 1480
rect 6908 140 6984 1480
rect 7188 140 7264 1480
rect 7468 140 7544 1480
rect 7748 140 7824 1480
rect 8028 140 8104 1480
rect 8308 140 8384 1480
rect 8588 140 8664 1480
rect 8868 140 8944 1480
rect 9148 140 9224 1480
rect 9428 0 9504 1620
use RM1 XRES1A
transform 1 0 200 0 1 202
box 200 202 320 202
use RM1 XRES1B
transform 1 0 200 0 1 1342
box 200 1342 320 1342
use RM1 XRES2
transform 1 0 200 0 1 658
box 200 658 320 658
use RM1 XRES4
transform 1 0 200 0 1 1114
box 200 1114 320 1114
use RM1 XRES8
transform 1 0 200 0 1 886
box 200 886 320 886
use RM1 XRES16
transform 1 0 200 0 1 430
box 200 430 320 430
use cut_M2M5_1x2 
transform 1 0 9428 0 1 610
box 9428 610 9504 810
use cut_M1M4_1x2 
transform 1 0 2428 0 1 140
box 2428 140 2504 340
use cut_M1M4_1x2 
transform 1 0 7188 0 1 1280
box 7188 1280 7264 1480
use cut_M1M4_1x2 
transform 1 0 2708 0 1 596
box 2708 596 2784 796
use cut_M1M4_1x2 
transform 1 0 6908 0 1 596
box 6908 596 6984 796
use cut_M1M4_1x2 
transform 1 0 2148 0 1 1052
box 2148 1052 2224 1252
use cut_M1M4_1x2 
transform 1 0 2988 0 1 1052
box 2988 1052 3064 1252
use cut_M1M4_1x2 
transform 1 0 6628 0 1 1052
box 6628 1052 6704 1252
use cut_M1M4_1x2 
transform 1 0 7468 0 1 1052
box 7468 1052 7544 1252
use cut_M1M4_1x2 
transform 1 0 1588 0 1 824
box 1588 824 1664 1024
use cut_M1M4_1x2 
transform 1 0 1868 0 1 824
box 1868 824 1944 1024
use cut_M1M4_1x2 
transform 1 0 3268 0 1 824
box 3268 824 3344 1024
use cut_M1M4_1x2 
transform 1 0 3548 0 1 824
box 3548 824 3624 1024
use cut_M1M4_1x2 
transform 1 0 6068 0 1 824
box 6068 824 6144 1024
use cut_M1M4_1x2 
transform 1 0 6348 0 1 824
box 6348 824 6424 1024
use cut_M1M4_1x2 
transform 1 0 7748 0 1 824
box 7748 824 7824 1024
use cut_M1M4_1x2 
transform 1 0 8028 0 1 824
box 8028 824 8104 1024
use cut_M1M4_1x2 
transform 1 0 468 0 1 368
box 468 368 544 568
use cut_M1M4_1x2 
transform 1 0 748 0 1 368
box 748 368 824 568
use cut_M1M4_1x2 
transform 1 0 1028 0 1 368
box 1028 368 1104 568
use cut_M1M4_1x2 
transform 1 0 1308 0 1 368
box 1308 368 1384 568
use cut_M1M4_1x2 
transform 1 0 3828 0 1 368
box 3828 368 3904 568
use cut_M1M4_1x2 
transform 1 0 4108 0 1 368
box 4108 368 4184 568
use cut_M1M4_1x2 
transform 1 0 4388 0 1 368
box 4388 368 4464 568
use cut_M1M4_1x2 
transform 1 0 4668 0 1 368
box 4668 368 4744 568
use cut_M1M4_1x2 
transform 1 0 4948 0 1 368
box 4948 368 5024 568
use cut_M1M4_1x2 
transform 1 0 5228 0 1 368
box 5228 368 5304 568
use cut_M1M4_1x2 
transform 1 0 5508 0 1 368
box 5508 368 5584 568
use cut_M1M4_1x2 
transform 1 0 5788 0 1 368
box 5788 368 5864 568
use cut_M1M4_1x2 
transform 1 0 8308 0 1 368
box 8308 368 8384 568
use cut_M1M4_1x2 
transform 1 0 8588 0 1 368
box 8588 368 8664 568
use cut_M1M4_1x2 
transform 1 0 8868 0 1 368
box 8868 368 8944 568
use cut_M1M4_1x2 
transform 1 0 9148 0 1 368
box 9148 368 9224 568
<< labels >>
flabel m3 s 328 0 404 1620 0 FreeSans 400 0 0 0 CTOP
port 7 nsew
flabel m1 s 328 0 9428 76 0 FreeSans 400 0 0 0 AVSS
port 8 nsew
flabel locali s 0 202 200 278 0 FreeSans 400 0 0 0 C1A
port 1 nsew
flabel locali s 0 1342 200 1418 0 FreeSans 400 0 0 0 C1B
port 2 nsew
flabel locali s 0 658 200 734 0 FreeSans 400 0 0 0 C2
port 3 nsew
flabel locali s 0 1114 200 1190 0 FreeSans 400 0 0 0 C4
port 4 nsew
flabel locali s 0 886 200 962 0 FreeSans 400 0 0 0 C8
port 5 nsew
flabel locali s 0 430 200 506 0 FreeSans 400 0 0 0 C16
port 6 nsew
<< end >>
