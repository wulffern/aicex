magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 1280
<< locali >>
rect 800 210 968 270
rect 800 850 968 910
rect 968 210 1520 270
rect 968 850 1520 910
rect 968 210 1028 910
rect 370 130 430 1150
rect 1890 130 1950 1150
rect 770 210 830 430
rect 770 530 830 750
rect 770 850 830 1070
rect 1490 210 1550 430
rect 1490 530 1550 750
rect 1490 850 1550 1070
<< poly >>
rect 280 142 2040 178
rect 280 462 2040 498
rect 280 782 2040 818
rect 280 1102 2040 1138
<< m2 >>
rect 1520 50 1688 110
rect 1520 530 1688 590
rect 1520 1170 1688 1230
rect 1688 530 2140 590
rect 1688 50 1748 1238
<< m3 >>
rect 680 0 880 1280
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1160 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1160 1280
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL MP2
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use PCHDL MP3
transform 1 0 1160 0 1 960
box 1160 960 2320 1280
use cut_M3M4_2x2 
transform 1 0 2040 0 1 530
box 2040 530 2240 730
use cut_M1M3_2x1 
transform 1 0 1400 0 1 50
box 1400 50 1600 118
use cut_M1M3_2x1 
transform 1 0 1400 0 1 530
box 1400 530 1600 598
use cut_M1M3_2x1 
transform 1 0 1400 0 1 1170
box 1400 1170 1600 1238
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
use cut_M1M4_2x1 
transform 1 0 680 0 1 530
box 680 530 880 598
use cut_M1M4_2x1 
transform 1 0 680 0 1 690
box 680 690 880 758
use cut_M1M4_2x1 
transform 1 0 680 0 1 1170
box 680 1170 880 1238
<< labels >>
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 680 210 920 270 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel m3 s 2040 530 2240 730 0 FreeSans 400 0 0 0 VREF
port 3 nsew
flabel m3 s 680 0 880 1280 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
<< end >>
