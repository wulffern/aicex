magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 1260 1760
<< locali >>
rect 402 146 462 1614
rect -108 132 108 220
rect 756 1642 972 1702
rect 324 146 540 206
rect 756 58 972 118
use SUNTR_NCHDL M0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_NCHDL M1
transform 1 0 0 0 1 176
box 0 176 1260 528
use SUNTR_NCHDL M2
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTR_NCHDL M3
transform 1 0 0 0 1 528
box 0 528 1260 880
use SUNTR_NCHDL M4
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNTR_NCHDL M5
transform 1 0 0 0 1 880
box 0 880 1260 1232
use SUNTR_NCHDL M6
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNTR_NCHDL M7
transform 1 0 0 0 1 1232
box 0 1232 1260 1584
use SUNTR_NCHDL M8
transform 1 0 0 0 1 1408
box 0 1408 1260 1760
<< labels >>
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 756 1642 972 1702 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 756 58 972 118 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
