magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 2360 4140
<< locali >>
rect 0 0 2360 112
rect 0 0 2360 112
rect 0 0 112 4140
rect 0 4028 2360 4140
rect 2248 0 2360 4140
rect 0 0 2360 112
rect 1450 3390 1774 3610
rect 586 3390 910 3610
<< ptapc >>
rect 20 0 100 80
rect 100 0 180 80
rect 180 0 260 80
rect 260 0 340 80
rect 340 0 420 80
rect 420 0 500 80
rect 500 0 580 80
rect 580 0 660 80
rect 660 0 740 80
rect 740 0 820 80
rect 820 0 900 80
rect 900 0 980 80
rect 980 0 1060 80
rect 1060 0 1140 80
rect 1140 0 1220 80
rect 1220 0 1300 80
rect 1300 0 1380 80
rect 1380 0 1460 80
rect 1460 0 1540 80
rect 1540 0 1620 80
rect 1620 0 1700 80
rect 1700 0 1780 80
rect 1780 0 1860 80
rect 1860 0 1940 80
rect 1940 0 2020 80
rect 2020 0 2100 80
rect 2100 0 2180 80
rect 2180 0 2260 80
rect 2260 0 2340 80
rect 0 30 80 110
rect 0 110 80 190
rect 0 190 80 270
rect 0 270 80 350
rect 0 350 80 430
rect 0 430 80 510
rect 0 510 80 590
rect 0 590 80 670
rect 0 670 80 750
rect 0 750 80 830
rect 0 830 80 910
rect 0 910 80 990
rect 0 990 80 1070
rect 0 1070 80 1150
rect 0 1150 80 1230
rect 0 1230 80 1310
rect 0 1310 80 1390
rect 0 1390 80 1470
rect 0 1470 80 1550
rect 0 1550 80 1630
rect 0 1630 80 1710
rect 0 1710 80 1790
rect 0 1790 80 1870
rect 0 1870 80 1950
rect 0 1950 80 2030
rect 0 2030 80 2110
rect 0 2110 80 2190
rect 0 2190 80 2270
rect 0 2270 80 2350
rect 0 2350 80 2430
rect 0 2430 80 2510
rect 0 2510 80 2590
rect 0 2590 80 2670
rect 0 2670 80 2750
rect 0 2750 80 2830
rect 0 2830 80 2910
rect 0 2910 80 2990
rect 0 2990 80 3070
rect 0 3070 80 3150
rect 0 3150 80 3230
rect 0 3230 80 3310
rect 0 3310 80 3390
rect 0 3390 80 3470
rect 0 3470 80 3550
rect 0 3550 80 3630
rect 0 3630 80 3710
rect 0 3710 80 3790
rect 0 3790 80 3870
rect 0 3870 80 3950
rect 0 3950 80 4030
rect 0 4030 80 4110
rect 20 4028 100 4108
rect 100 4028 180 4108
rect 180 4028 260 4108
rect 260 4028 340 4108
rect 340 4028 420 4108
rect 420 4028 500 4108
rect 500 4028 580 4108
rect 580 4028 660 4108
rect 660 4028 740 4108
rect 740 4028 820 4108
rect 820 4028 900 4108
rect 900 4028 980 4108
rect 980 4028 1060 4108
rect 1060 4028 1140 4108
rect 1140 4028 1220 4108
rect 1220 4028 1300 4108
rect 1300 4028 1380 4108
rect 1380 4028 1460 4108
rect 1460 4028 1540 4108
rect 1540 4028 1620 4108
rect 1620 4028 1700 4108
rect 1700 4028 1780 4108
rect 1780 4028 1860 4108
rect 1860 4028 1940 4108
rect 1940 4028 2020 4108
rect 2020 4028 2100 4108
rect 2100 4028 2180 4108
rect 2180 4028 2260 4108
rect 2260 4028 2340 4108
rect 2248 30 2328 110
rect 2248 110 2328 190
rect 2248 190 2328 270
rect 2248 270 2328 350
rect 2248 350 2328 430
rect 2248 430 2328 510
rect 2248 510 2328 590
rect 2248 590 2328 670
rect 2248 670 2328 750
rect 2248 750 2328 830
rect 2248 830 2328 910
rect 2248 910 2328 990
rect 2248 990 2328 1070
rect 2248 1070 2328 1150
rect 2248 1150 2328 1230
rect 2248 1230 2328 1310
rect 2248 1310 2328 1390
rect 2248 1390 2328 1470
rect 2248 1470 2328 1550
rect 2248 1550 2328 1630
rect 2248 1630 2328 1710
rect 2248 1710 2328 1790
rect 2248 1790 2328 1870
rect 2248 1870 2328 1950
rect 2248 1950 2328 2030
rect 2248 2030 2328 2110
rect 2248 2110 2328 2190
rect 2248 2190 2328 2270
rect 2248 2270 2328 2350
rect 2248 2350 2328 2430
rect 2248 2430 2328 2510
rect 2248 2510 2328 2590
rect 2248 2590 2328 2670
rect 2248 2670 2328 2750
rect 2248 2750 2328 2830
rect 2248 2830 2328 2910
rect 2248 2910 2328 2990
rect 2248 2990 2328 3070
rect 2248 3070 2328 3150
rect 2248 3150 2328 3230
rect 2248 3230 2328 3310
rect 2248 3310 2328 3390
rect 2248 3390 2328 3470
rect 2248 3470 2328 3550
rect 2248 3550 2328 3630
rect 2248 3630 2328 3710
rect 2248 3710 2328 3790
rect 2248 3790 2328 3870
rect 2248 3870 2328 3950
rect 2248 3950 2328 4030
rect 2248 4030 2328 4110
<< ptap >>
rect 0 0 2360 112
rect 0 0 112 4140
rect 0 4028 2360 4140
rect 2248 0 2360 4140
use SUNTR_RES25 XA1
transform 1 0 640 0 1 640
box 640 640 1720 3500
<< labels >>
flabel locali s 0 0 2360 112 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 1450 3390 1774 3610 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 586 3390 910 3610 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
