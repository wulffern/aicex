
*-------------------------------------------------------------
* SUNTR_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLR D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLCM D G S B
XM0 N0 G S B SUNTR_NCHDL
XM1 N1 G N0 B SUNTR_NCHDL
XM2 N2 G N1 B SUNTR_NCHDL
XM3 N3 G N2 B SUNTR_NCHDL
XM4 N4 G N3 B SUNTR_NCHDL
XM5 N5 G N4 B SUNTR_NCHDL
XM6 N6 G N5 B SUNTR_NCHDL
XM7 N7 G N6 B SUNTR_NCHDL
XM8 D G N7 B SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLCM D G S B
XM0 N0 G S B SUNTR_PCHDL
XM7 D G N0 B SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLA D G S B
XM0 D G S B SUNTR_NCHDL
XM1 S G D B SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLA D G S B
XM0 D G S B SUNTR_PCHDL
XM1 S G D B SUNTR_PCHDL
XM2 D G S B SUNTR_PCHDL
XM3 S G D B SUNTR_PCHDL
XM4 D G S B SUNTR_PCHDL
XM5 S G D B SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLCM2 D G S B
XM0 D G S B SUNTR_NCHDLCM
XM1 S G D B SUNTR_NCHDLCM
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLCM2 D G S B
XM0 D G S B SUNTR_PCHDLCM
XM1 S G D B SUNTR_PCHDLCM
.ENDS

*-------------------------------------------------------------
* SUNTR_CPCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_CPCHDLCM2 D G CG S CS B
XM0 CS G S B SUNTR_PCHDLCM2
XM1 D CG CS B SUNTR_PCHDLA
.ENDS

*-------------------------------------------------------------
* SUNTR_CNCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_CNCHDLCM2 D G CG S CS B
XM0 CS G S B SUNTR_NCHDLCM2
XM1 D CG CS B SUNTR_NCHDLA
.ENDS

*-------------------------------------------------------------
* SUNTR_TAPCELLB_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTR_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_TIEH_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TIEH_CV Y AVDD AVSS
XMN0 A A AVSS AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_TIEL_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TIEL_CV Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMP0 A A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX1_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX2_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX4_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
XMP2 Y A AVDD AVDD SUNTR_PCHDL
XMP3 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX8_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMN4 Y A AVSS AVSS SUNTR_NCHDL
XMN5 AVSS A Y AVSS SUNTR_NCHDL
XMN6 Y A AVSS AVSS SUNTR_NCHDL
XMN7 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
XMP2 Y A AVDD AVDD SUNTR_PCHDL
XMP3 AVDD A Y AVDD SUNTR_PCHDL
XMP4 Y A AVDD AVDD SUNTR_PCHDL
XMP5 AVDD A Y AVDD SUNTR_PCHDL
XMP6 Y A AVDD AVDD SUNTR_PCHDL
XMP7 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_BFX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_BFX1_CV A Y AVDD AVSS
XMN0 AVSS A B AVSS SUNTR_NCHDL
XMN1 Y B AVSS AVSS SUNTR_NCHDL
XMP0 AVDD A B AVDD SUNTR_PCHDL
XMP1 Y B AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NRX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NRX1_CV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS B Y AVSS SUNTR_NCHDL
XMP0 N1 A AVDD AVDD SUNTR_PCHDL
XMP1 Y B N1 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NDX1_CV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y B N1 AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD B Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_ORX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ORX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NRX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ORX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ORX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NRX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ORX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ORX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NRX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX8_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_IVTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVTRIX1_CV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y C N1 AVSS SUNTR_NCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NDTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NDTRIX1_CV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS SUNTR_NCHDL
XMN0 N2 A N1 AVSS SUNTR_NCHDL
XMN1 Y C N2 AVSS SUNTR_NCHDL
XMP2 AVDD RN N2 AVDD SUNTR_PCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NRTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NRTRIX1_CV A C CN B Y AVDD AVSS
XMN2 N1 B AVSS AVSS SUNTR_NCHDL
XMN0 AVSS A N1 AVSS SUNTR_NCHDL
XMN1 N1 C Y AVSS SUNTR_NCHDL
XMP2 N2 B AVDD AVDD SUNTR_PCHDL
XMP0 AVDD A N2 AVDD SUNTR_PCHDL
XMP1 N2 CN Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_DFRNQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS SUNTR_TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS SUNTR_NDX1_CV
XA2 CKN CKB AVDD AVSS SUNTR_IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS SUNTR_IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS SUNTR_IVTRIX1_CV
XA5 A0 A1 AVDD AVSS SUNTR_IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS SUNTR_IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS SUNTR_NDTRIX1_CV
XA8 QN Q AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_SCX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SCX1_CV A Y AVDD AVSS
XA2 N1 A AVSS AVSS SUNTR_NCHDL
XA3 SCO A N1 AVSS SUNTR_NCHDL
XA4a AVDD SCO N1 AVSS SUNTR_NCHDL
XA4b AVDD SCO N1 AVSS SUNTR_NCHDL
XA5 Y SCO AVSS AVSS SUNTR_NCHDL
XB0 N2 A AVDD AVDD SUNTR_PCHDL
XB1 SCO A N2 AVDD SUNTR_PCHDL
XB3a N2 SCO AVSS AVDD SUNTR_PCHDL
XB3b N2 SCO AVSS AVDD SUNTR_PCHDL
XB4 Y SCO AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_SWX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SWX2_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A VREF AVDD SUNTR_PCHDL
XMP1 VREF A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_SWX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SWX4_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A VREF AVDD SUNTR_PCHDL
XMP1 VREF A Y AVDD SUNTR_PCHDL
XMP2 Y A VREF AVDD SUNTR_PCHDL
XMP3 VREF A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_TGPD_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TGPD_CV C A B AVDD AVSS
XMN0 AVSS C CN AVSS SUNTR_NCHDL
XMN1 B C AVSS AVSS SUNTR_NCHDL
XMN2 A CN B AVSS SUNTR_NCHDL
XMP0 AVDD C CN AVDD SUNTR_PCHDL
XMP1_DMY B AVDD AVDD AVDD SUNTR_PCHDL
XMP2 A C B AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_DFTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFTRIX1_CV D CK C CN Y AVDD AVSS
XA3 AVDD AVSS SUNTR_TAPCELLB_CV
XA2 D CK C NC QN AVDD AVSS SUNTR_DFRNQNX1_CV
XA0 QN C CN Y AVDD AVSS SUNTR_IVTRIX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_RG12TRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RG12TRIX1_CV D<11> D<10> D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> CK C CN Y<11> Y<10> Y<9> Y<8> Y<7> Y<6> Y<5> Y<4> Y<3> Y<2> Y<1> Y<0> AVDD AVSS
XA0 D<11> CK C CN Y<11> AVDD AVSS SUNTR_DFTRIX1_CV
XB1 D<10> CK C CN Y<10> AVDD AVSS SUNTR_DFTRIX1_CV
XC2 D<9> CK C CN Y<9> AVDD AVSS SUNTR_DFTRIX1_CV
XD3 D<8> CK C CN Y<8> AVDD AVSS SUNTR_DFTRIX1_CV
XE4 D<7> CK C CN Y<7> AVDD AVSS SUNTR_DFTRIX1_CV
XF5 D<6> CK C CN Y<6> AVDD AVSS SUNTR_DFTRIX1_CV
XG6 D<5> CK C CN Y<5> AVDD AVSS SUNTR_DFTRIX1_CV
XH7 D<4> CK C CN Y<4> AVDD AVSS SUNTR_DFTRIX1_CV
XI8 D<3> CK C CN Y<3> AVDD AVSS SUNTR_DFTRIX1_CV
XJ9 D<2> CK C CN Y<2> AVDD AVSS SUNTR_DFTRIX1_CV
XK10 D<1> CK C CN Y<1> AVDD AVSS SUNTR_DFTRIX1_CV
XL11 D<0> CK C CN Y<0> AVDD AVSS SUNTR_DFTRIX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_SUN_TR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SUN_TR AVDD AVSS
XA0 AVDD AVSS SUNTR_TAPCELLB_CV
XA1 Y1 AVDD AVSS SUNTR_TIEH_CV
XA2 Y2 AVDD AVSS SUNTR_TIEL_CV
XB0 AVDD AVSS SUNTR_TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS SUNTR_IVX1_CV
XB4 A4 Y4 AVDD AVSS SUNTR_IVX2_CV
XB5 A5 Y5 AVDD AVSS SUNTR_IVX4_CV
XB6 A6 Y6 AVDD AVSS SUNTR_IVX8_CV
XC0 AVDD AVSS SUNTR_TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS SUNTR_BFX1_CV
XD0 AVDD AVSS SUNTR_TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS SUNTR_NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS SUNTR_NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS SUNTR_ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS SUNTR_ANX1_CV
XE0 AVDD AVSS SUNTR_TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SUNTR_SCX1_CV
XF0 AVDD AVSS SUNTR_TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SUNTR_SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SUNTR_SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS SUNTR_TGPD_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTRB_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTRB_NCHDLR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NCHDLR D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTRB_TIEH_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_TIEH_CV Y BULKP BULKN AVDD AVSS
XMN0 A A AVSS BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_TIEL_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_TIEL_CV Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMP0 A A AVDD BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_IVX1_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_IVX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_IVX2_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMN1 AVSS A Y BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
XMP1 AVDD A Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_IVX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_IVX4_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMN1 AVSS A Y BULKN SUNTRB_NCHDL
XMN2 Y A AVSS BULKN SUNTRB_NCHDL
XMN3 AVSS A Y BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
XMP1 AVDD A Y BULKP SUNTRB_PCHDL
XMP2 Y A AVDD BULKP SUNTRB_PCHDL
XMP3 AVDD A Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_IVX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_IVX8_CV A Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMN1 AVSS A Y BULKN SUNTRB_NCHDL
XMN2 Y A AVSS BULKN SUNTRB_NCHDL
XMN3 AVSS A Y BULKN SUNTRB_NCHDL
XMN4 Y A AVSS BULKN SUNTRB_NCHDL
XMN5 AVSS A Y BULKN SUNTRB_NCHDL
XMN6 Y A AVSS BULKN SUNTRB_NCHDL
XMN7 AVSS A Y BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
XMP1 AVDD A Y BULKP SUNTRB_PCHDL
XMP2 Y A AVDD BULKP SUNTRB_PCHDL
XMP3 AVDD A Y BULKP SUNTRB_PCHDL
XMP4 Y A AVDD BULKP SUNTRB_PCHDL
XMP5 AVDD A Y BULKP SUNTRB_PCHDL
XMP6 Y A AVDD BULKP SUNTRB_PCHDL
XMP7 AVDD A Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_BFX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_BFX1_CV A Y BULKP BULKN AVDD AVSS
XMN0 AVSS A B BULKN SUNTRB_NCHDL
XMN1 Y B AVSS BULKN SUNTRB_NCHDL
XMP0 AVDD A B BULKP SUNTRB_PCHDL
XMP1 Y B AVDD BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_NRX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NRX1_CV A B Y BULKP BULKN AVDD AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMN1 AVSS B Y BULKN SUNTRB_NCHDL
XMP0 N1 A AVDD BULKP SUNTRB_PCHDL
XMP1 Y B N1 BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NDX1_CV A B Y BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNTRB_NCHDL
XMN1 Y B N1 BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
XMP1 AVDD B Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_ORX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ORX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_ORX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ORX2_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX2_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_ORX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ORX4_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NRX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX4_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_ANX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ANX1_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_ANX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ANX2_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX2_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_ANX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ANX4_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX4_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_ANX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_ANX8_CV A B Y BULKP BULKN AVDD AVSS
XA1 A B YN BULKP BULKN AVDD AVSS SUNTRB_NDX1_CV
XA2 YN Y BULKP BULKN AVDD AVSS SUNTRB_IVX8_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_IVTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_IVTRIX1_CV A C CN Y BULKP BULKN AVDD AVSS
XMN0 N1 A AVSS BULKN SUNTRB_NCHDL
XMN1 Y C N1 BULKN SUNTRB_NCHDL
XMP0 N2 A AVDD BULKP SUNTRB_PCHDL
XMP1 Y CN N2 BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_NDTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_NDTRIX1_CV A C CN RN Y BULKP BULKN AVDD AVSS
XMN2 N1 RN AVSS BULKN SUNTRB_NCHDL
XMN0 N2 A N1 BULKN SUNTRB_NCHDL
XMN1 Y C N2 BULKN SUNTRB_NCHDL
XMP2 AVDD RN N2 BULKP SUNTRB_PCHDL
XMP0 N2 A AVDD BULKP SUNTRB_PCHDL
XMP1 Y CN N2 BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_DFRNQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_DFRNQNX1_CV D CK RN Q QN BULKP BULKN AVDD AVSS
XA0 BULKP BULKN SUNTRB_TAPCELLB_CV
XA1 CK RN CKN BULKP BULKN AVDD AVSS SUNTRB_NDX1_CV
XA2 CKN CKB BULKP BULKN AVDD AVSS SUNTRB_IVX1_CV
XA3 D CKN CKB A0 BULKP BULKN AVDD AVSS SUNTRB_IVTRIX1_CV
XA4 A1 CKB CKN A0 BULKP BULKN AVDD AVSS SUNTRB_IVTRIX1_CV
XA5 A0 A1 BULKP BULKN AVDD AVSS SUNTRB_IVX1_CV
XA6 A1 CKB CKN QN BULKP BULKN AVDD AVSS SUNTRB_IVTRIX1_CV
XA7 Q CKN CKB RN QN BULKP BULKN AVDD AVSS SUNTRB_NDTRIX1_CV
XA8 QN Q BULKP BULKN AVDD AVSS SUNTRB_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTRB_SCX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_SCX1_CV A Y BULKP BULKN AVDD AVSS
XA2 N1 A AVSS BULKN SUNTRB_NCHDL
XA3 SCO A N1 BULKN SUNTRB_NCHDL
XA4a AVDD SCO N1 BULKN SUNTRB_NCHDL
XA4b AVDD SCO N1 BULKN SUNTRB_NCHDL
XA5 Y SCO AVSS BULKN SUNTRB_NCHDL
XB0 N2 A AVDD BULKP SUNTRB_PCHDL
XB1 SCO A N2 BULKP SUNTRB_PCHDL
XB3a N2 SCO AVSS BULKP SUNTRB_PCHDL
XB3b N2 SCO AVSS BULKP SUNTRB_PCHDL
XB4 Y SCO AVDD AVSS SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_SWX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_SWX2_CV A Y VREF AVSS BULKP BULKN
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMN1 AVSS A Y BULKN SUNTRB_NCHDL
XMP0 Y A VREF BULKP SUNTRB_PCHDL
XMP1 VREF A Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_SWX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_SWX4_CV A Y VREF AVSS BULKP BULKN
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMN1 AVSS A Y BULKN SUNTRB_NCHDL
XMN2 Y A AVSS BULKN SUNTRB_NCHDL
XMN3 AVSS A Y BULKN SUNTRB_NCHDL
XMP0 Y A VREF BULKP SUNTRB_PCHDL
XMP1 VREF A Y BULKP SUNTRB_PCHDL
XMP2 Y A VREF BULKP SUNTRB_PCHDL
XMP3 VREF A Y BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_TGPD_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_TGPD_CV C A B BULKP BULKN AVDD AVSS
XMN0 AVSS C CN BULKN SUNTRB_NCHDL
XMN1 B C AVSS BULKN SUNTRB_NCHDL
XMN2 A CN B BULKN SUNTRB_NCHDL
XMP0 AVDD C CN BULKP SUNTRB_PCHDL
XMP1_DMY B AVDD AVDD BULKP SUNTRB_PCHDL
XMP2 A C B BULKP SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_TAPCELLB_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTRB_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTRB_TAPCELLBAVSS_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTRB_TAPCELLBAVSS_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTRB_NCHDL
XMP1 NC1 NC1 NC1 AVDD SUNTRB_PCHDL
.ENDS

*-------------------------------------------------------------
* SUN_PLL_LSCORE <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_LSCORE A AN YN Y AVDD AVSS
xb1_0 Y AN AVSS AVSS SUNTR_NCHDL
xb1_1 Y AN AVSS AVSS SUNTR_NCHDL
xb2_0 YN A AVSS AVSS SUNTR_NCHDL
xb2_1 YN A AVSS AVSS SUNTR_NCHDL
xc1a net2 YN AVDD AVDD SUNTR_PCHDL
xc1b Y YN net2 AVDD SUNTR_PCHDL
xc2a net1 Y AVDD AVDD SUNTR_PCHDL
xc2b YN Y net1 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUN_PLL_ROSC <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUN_PLL_ROSC PWRUP_1V8 VDD_ROSC AVSS VDD_1V8 CK
xa3 N_2 N_1 CKUP NC1 VDD_1V8 AVSS SUN_PLL_LSCORE
xa4 CKUP CK VDD_1V8 AVSS SUNTR_IVX1_CV
xa5 VDD_1V8 AVSS SUNTR_TAPCELLB_CV
xb1 PWRUP_1V8 N_0 NI VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_NDX1_CV
xb2_0 NI N_7 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_1 N_7 N_6 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_2 N_6 N_5 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_3 N_5 N_4 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_4 N_4 N_3 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_5 N_3 N_2 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_6 N_2 N_1 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_7 N_1 N_0 VDD_1V8 AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb3 VDD_1V8 AVSS SUNTRB_TAPCELLBAVSS_CV
.ENDS
