magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 1600
<< locali >>
rect 720 210 858 270
rect 720 370 858 430
rect 720 690 858 750
rect 720 1010 858 1070
rect 858 210 918 1070
rect 1062 210 1260 270
rect 1062 370 1260 430
rect 1062 850 1260 910
rect 1062 1170 1260 1230
rect 1062 210 1122 1230
rect 330 130 390 510
rect 1620 770 1758 830
rect 1260 530 1758 590
rect 1620 1090 1758 1150
rect 1620 1410 1758 1470
rect 1758 530 1818 1470
rect 162 770 360 830
rect 162 530 720 590
rect 162 1090 360 1150
rect 162 1410 360 1470
rect 162 530 222 1470
rect 522 850 720 910
rect 522 1170 720 1230
rect 522 850 582 1230
rect 720 1490 858 1550
rect 858 1490 1260 1550
rect 858 1490 918 1550
rect 720 1170 858 1230
rect 858 1330 1260 1390
rect 858 1170 918 1390
rect 1260 690 1398 750
rect 1260 1010 1398 1070
rect 1398 690 1458 1070
<< m1 >>
rect 720 1330 858 1390
rect 858 1010 1260 1070
rect 858 1010 918 1398
rect 720 530 858 590
rect 858 530 1260 590
rect 858 530 918 598
<< poly >>
rect 270 142 1710 178
rect 270 462 1710 498
<< m3 >>
rect 1170 0 1354 1600
rect 630 0 814 1600
use NCHDL XA2
transform 1 0 0 0 1 0
box 0 0 990 320
use NCHDL XA3
transform 1 0 0 0 1 320
box 0 320 990 640
use NCHDL XA4a
transform 1 0 0 0 1 640
box 0 640 990 960
use NCHDL XA4b
transform 1 0 0 0 1 960
box 0 960 990 1280
use NCHDL XA5
transform 1 0 0 0 1 1280
box 0 1280 990 1600
use PCHDL XB0
transform 1 0 990 0 1 0
box 990 0 1980 320
use PCHDL XB1
transform 1 0 990 0 1 320
box 990 320 1980 640
use PCHDL XB3a
transform 1 0 990 0 1 640
box 990 640 1980 960
use PCHDL XB3b
transform 1 0 990 0 1 960
box 990 960 1980 1280
use PCHDL XB4
transform 1 0 990 0 1 1280
box 990 1280 1980 1600
use cut_M1M2_2x1 
transform 1 0 630 0 1 1330
box 630 1330 814 1398
use cut_M1M2_2x1 
transform 1 0 1170 0 1 1010
box 1170 1010 1354 1078
use cut_M1M2_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M2_2x1 
transform 1 0 1170 0 1 530
box 1170 530 1354 598
use cut_M1M4_2x1 
transform 1 0 1170 0 1 50
box 1170 50 1354 118
use cut_M1M4_2x1 
transform 1 0 1170 0 1 1330
box 1170 1330 1354 1398
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 1330
box 630 1330 814 1398
<< labels >>
flabel locali s 270 130 450 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 630 1490 810 1550 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel m3 s 1170 0 1354 1600 0 FreeSans 400 0 0 0 AVDD
port 3 nsew
flabel m3 s 630 0 814 1600 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
<< end >>
