magic
tech sky130A
magscale 1 2
timestamp 1658699483
<< checkpaint >>
rect 0 0 184 68
<< locali >>
rect 0 0 184 68
<< m1 >>
rect 0 0 184 68
<< viali >>
rect 12 6 172 62
<< labels >>
<< end >>
