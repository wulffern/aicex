magic
tech sky130A
magscale 1 2
timestamp 1661983200
<< checkpaint >>
rect 0 0 40696 26808
<< locali >>
rect 40396 0 40696 26808
rect 0 0 40696 300
rect 0 26508 40696 26808
rect 0 0 300 26808
rect 40396 0 40696 26808
rect 300 636 460 748
rect 300 5048 460 5160
rect 300 9460 460 9572
rect 300 13872 460 13984
rect 300 18284 460 18396
rect 5380 21706 5956 21926
rect 1060 4058 1636 4278
<< m3 >>
rect 23264 0 23480 484
rect 40132 404 40472 480
rect 40132 1364 40472 1440
rect 40132 2324 40472 2400
rect 40132 3284 40472 3360
rect 40132 4244 40472 4320
rect 40132 5204 40472 5280
rect 40132 6164 40472 6240
rect 40132 7124 40472 7200
rect 40132 8084 40472 8160
rect 40132 9044 40472 9120
rect 40132 10004 40472 10080
rect 40132 10964 40472 11040
rect 40132 11924 40472 12000
rect 40132 12884 40472 12960
rect 40132 13844 40472 13920
rect 40132 14804 40472 14880
rect 40132 15764 40472 15840
rect 40132 16724 40472 16800
rect 40132 17684 40472 17760
rect 40132 18644 40472 18720
rect 40132 19604 40472 19680
rect 40132 20564 40472 20640
rect 40132 21524 40472 21600
rect 40132 22484 40472 22560
rect 40132 23444 40472 23520
rect 40132 24404 40472 24480
rect 40132 25364 40472 25440
<< m1 >>
rect 1152 8470 1364 8530
rect 1364 4058 5472 4118
rect 1364 4058 1424 8538
rect 1152 17294 1508 17354
rect 1508 12882 5472 12942
rect 1508 12882 1568 17362
rect 5472 21706 5624 21766
rect 5624 4084 6712 4144
rect 5624 5044 6712 5104
rect 5624 6004 6712 6064
rect 5624 6964 6712 7024
rect 5624 7924 6712 7984
rect 5624 8884 6712 8944
rect 5624 9844 6712 9904
rect 5624 10804 6712 10864
rect 5624 11764 6712 11824
rect 5624 12724 6712 12784
rect 5624 13684 6712 13744
rect 5624 14644 6712 14704
rect 5624 15604 6712 15664
rect 5624 16564 6712 16624
rect 5624 17524 6712 17584
rect 5624 18484 6712 18544
rect 5624 19444 6712 19504
rect 5624 20404 6712 20464
rect 5624 21364 6712 21424
rect 5624 22324 6712 22384
rect 5624 23284 6712 23344
rect 5624 24244 6712 24304
rect 5624 25204 6712 25264
rect 5624 26164 6712 26224
rect 5624 4084 5684 26240
<< m2 >>
rect 1160 12882 1388 12958
rect 1388 8470 5480 8546
rect 1388 8470 1464 12958
rect 1160 21706 1676 21782
rect 1676 17294 5480 17370
rect 1676 17294 1752 21782
rect 1160 4058 1324 4134
rect 1324 1204 6712 1280
rect 1324 2164 6712 2240
rect 1324 3124 6712 3200
rect 1324 1204 1400 4134
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa10
transform 1 0 444 0 1 620
box 444 620 6572 4856
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa20
transform 1 0 444 0 1 5032
box 444 5032 6572 9268
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa30
transform 1 0 444 0 1 9444
box 444 9444 6572 13680
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa40
transform 1 0 444 0 1 13856
box 444 13856 6572 18092
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa50
transform 1 0 444 0 1 18268
box 444 18268 6572 22504
use CAP_LPF xb10
transform -1 0 40252 0 1 444
box 40252 444 73932 1404
use CAP_LPF xb20
transform -1 0 40252 0 1 1404
box 40252 1404 73932 2364
use CAP_LPF xb21
transform -1 0 40252 0 1 2364
box 40252 2364 73932 3324
use CAP_LPF xb30
transform -1 0 40252 0 1 3324
box 40252 3324 73932 4284
use CAP_LPF xb31
transform -1 0 40252 0 1 4284
box 40252 4284 73932 5244
use CAP_LPF xb32
transform -1 0 40252 0 1 5244
box 40252 5244 73932 6204
use CAP_LPF xb33
transform -1 0 40252 0 1 6204
box 40252 6204 73932 7164
use CAP_LPF xb34
transform -1 0 40252 0 1 7164
box 40252 7164 73932 8124
use CAP_LPF xb35
transform -1 0 40252 0 1 8124
box 40252 8124 73932 9084
use CAP_LPF xb36
transform -1 0 40252 0 1 9084
box 40252 9084 73932 10044
use CAP_LPF xb37
transform -1 0 40252 0 1 10044
box 40252 10044 73932 11004
use CAP_LPF xb38
transform -1 0 40252 0 1 11004
box 40252 11004 73932 11964
use CAP_LPF xb39
transform -1 0 40252 0 1 11964
box 40252 11964 73932 12924
use CAP_LPF xb310
transform -1 0 40252 0 1 12924
box 40252 12924 73932 13884
use CAP_LPF xb311
transform -1 0 40252 0 1 13884
box 40252 13884 73932 14844
use CAP_LPF xb312
transform -1 0 40252 0 1 14844
box 40252 14844 73932 15804
use CAP_LPF xb313
transform -1 0 40252 0 1 15804
box 40252 15804 73932 16764
use CAP_LPF xb314
transform -1 0 40252 0 1 16764
box 40252 16764 73932 17724
use CAP_LPF xb315
transform -1 0 40252 0 1 17724
box 40252 17724 73932 18684
use CAP_LPF xb316
transform -1 0 40252 0 1 18684
box 40252 18684 73932 19644
use CAP_LPF xb317
transform -1 0 40252 0 1 19644
box 40252 19644 73932 20604
use CAP_LPF xb318
transform -1 0 40252 0 1 20604
box 40252 20604 73932 21564
use CAP_LPF xb319
transform -1 0 40252 0 1 21564
box 40252 21564 73932 22524
use CAP_LPF xb320
transform -1 0 40252 0 1 22524
box 40252 22524 73932 23484
use CAP_LPF xb321
transform -1 0 40252 0 1 23484
box 40252 23484 73932 24444
use CAP_LPF xb322
transform -1 0 40252 0 1 24444
box 40252 24444 73932 25404
use CAP_LPF xb323
transform -1 0 40252 0 1 25404
box 40252 25404 73932 26364
use cut_M1M4_2x1 
transform 1 0 23272 0 1 0
box 23272 0 23472 76
use cut_M1M2_2x1 
transform 1 0 1060 0 1 8470
box 1060 8470 1244 8538
use cut_M1M2_2x1 
transform 1 0 5380 0 1 4058
box 5380 4058 5564 4126
use cut_M1M3_2x1 
transform 1 0 1060 0 1 12882
box 1060 12882 1260 12958
use cut_M1M3_2x1 
transform 1 0 5380 0 1 8470
box 5380 8470 5580 8546
use cut_M1M2_2x1 
transform 1 0 1060 0 1 17294
box 1060 17294 1244 17362
use cut_M1M2_2x1 
transform 1 0 5380 0 1 12882
box 5380 12882 5564 12950
use cut_M1M3_2x1 
transform 1 0 1060 0 1 21706
box 1060 21706 1260 21782
use cut_M1M3_2x1 
transform 1 0 5380 0 1 17294
box 5380 17294 5580 17370
use cut_M1M2_2x1 
transform 1 0 5380 0 1 21706
box 5380 21706 5564 21774
use cut_M2M4_2x1 
transform 1 0 6612 0 1 4084
box 6612 4084 6812 4160
use cut_M2M4_2x1 
transform 1 0 6612 0 1 5044
box 6612 5044 6812 5120
use cut_M2M4_2x1 
transform 1 0 6612 0 1 6004
box 6612 6004 6812 6080
use cut_M2M4_2x1 
transform 1 0 6612 0 1 6964
box 6612 6964 6812 7040
use cut_M2M4_2x1 
transform 1 0 6612 0 1 7924
box 6612 7924 6812 8000
use cut_M2M4_2x1 
transform 1 0 6612 0 1 8884
box 6612 8884 6812 8960
use cut_M2M4_2x1 
transform 1 0 6612 0 1 9844
box 6612 9844 6812 9920
use cut_M2M4_2x1 
transform 1 0 6612 0 1 10804
box 6612 10804 6812 10880
use cut_M2M4_2x1 
transform 1 0 6612 0 1 11764
box 6612 11764 6812 11840
use cut_M2M4_2x1 
transform 1 0 6612 0 1 12724
box 6612 12724 6812 12800
use cut_M2M4_2x1 
transform 1 0 6612 0 1 13684
box 6612 13684 6812 13760
use cut_M2M4_2x1 
transform 1 0 6612 0 1 14644
box 6612 14644 6812 14720
use cut_M2M4_2x1 
transform 1 0 6612 0 1 15604
box 6612 15604 6812 15680
use cut_M2M4_2x1 
transform 1 0 6612 0 1 16564
box 6612 16564 6812 16640
use cut_M2M4_2x1 
transform 1 0 6612 0 1 17524
box 6612 17524 6812 17600
use cut_M2M4_2x1 
transform 1 0 6612 0 1 18484
box 6612 18484 6812 18560
use cut_M2M4_2x1 
transform 1 0 6612 0 1 19444
box 6612 19444 6812 19520
use cut_M2M4_2x1 
transform 1 0 6612 0 1 20404
box 6612 20404 6812 20480
use cut_M2M4_2x1 
transform 1 0 6612 0 1 21364
box 6612 21364 6812 21440
use cut_M2M4_2x1 
transform 1 0 6612 0 1 22324
box 6612 22324 6812 22400
use cut_M2M4_2x1 
transform 1 0 6612 0 1 23284
box 6612 23284 6812 23360
use cut_M2M4_2x1 
transform 1 0 6612 0 1 24244
box 6612 24244 6812 24320
use cut_M2M4_2x1 
transform 1 0 6612 0 1 25204
box 6612 25204 6812 25280
use cut_M2M4_2x1 
transform 1 0 6612 0 1 26164
box 6612 26164 6812 26240
use cut_M1M3_2x1 
transform 1 0 1060 0 1 4058
box 1060 4058 1260 4134
use cut_M3M4_2x1 
transform 1 0 6612 0 1 1204
box 6612 1204 6812 1280
use cut_M3M4_2x1 
transform 1 0 6612 0 1 2164
box 6612 2164 6812 2240
use cut_M3M4_2x1 
transform 1 0 6612 0 1 3124
box 6612 3124 6812 3200
use cut_M1M4_1x2 
transform 1 0 40396 0 1 0
box 40396 0 40472 200
use cut_M1M4_1x2 
transform 1 0 40396 0 1 404
box 40396 404 40472 604
use cut_M1M4_1x2 
transform 1 0 40396 0 1 1364
box 40396 1364 40472 1564
use cut_M1M4_1x2 
transform 1 0 40396 0 1 2324
box 40396 2324 40472 2524
use cut_M1M4_1x2 
transform 1 0 40396 0 1 3284
box 40396 3284 40472 3484
use cut_M1M4_1x2 
transform 1 0 40396 0 1 4244
box 40396 4244 40472 4444
use cut_M1M4_1x2 
transform 1 0 40396 0 1 5204
box 40396 5204 40472 5404
use cut_M1M4_1x2 
transform 1 0 40396 0 1 6164
box 40396 6164 40472 6364
use cut_M1M4_1x2 
transform 1 0 40396 0 1 7124
box 40396 7124 40472 7324
use cut_M1M4_1x2 
transform 1 0 40396 0 1 8084
box 40396 8084 40472 8284
use cut_M1M4_1x2 
transform 1 0 40396 0 1 9044
box 40396 9044 40472 9244
use cut_M1M4_1x2 
transform 1 0 40396 0 1 10004
box 40396 10004 40472 10204
use cut_M1M4_1x2 
transform 1 0 40396 0 1 10964
box 40396 10964 40472 11164
use cut_M1M4_1x2 
transform 1 0 40396 0 1 11924
box 40396 11924 40472 12124
use cut_M1M4_1x2 
transform 1 0 40396 0 1 12884
box 40396 12884 40472 13084
use cut_M1M4_1x2 
transform 1 0 40396 0 1 13844
box 40396 13844 40472 14044
use cut_M1M4_1x2 
transform 1 0 40396 0 1 14804
box 40396 14804 40472 15004
use cut_M1M4_1x2 
transform 1 0 40396 0 1 15764
box 40396 15764 40472 15964
use cut_M1M4_1x2 
transform 1 0 40396 0 1 16724
box 40396 16724 40472 16924
use cut_M1M4_1x2 
transform 1 0 40396 0 1 17684
box 40396 17684 40472 17884
use cut_M1M4_1x2 
transform 1 0 40396 0 1 18644
box 40396 18644 40472 18844
use cut_M1M4_1x2 
transform 1 0 40396 0 1 19604
box 40396 19604 40472 19804
use cut_M1M4_1x2 
transform 1 0 40396 0 1 20564
box 40396 20564 40472 20764
use cut_M1M4_1x2 
transform 1 0 40396 0 1 21524
box 40396 21524 40472 21724
use cut_M1M4_1x2 
transform 1 0 40396 0 1 22484
box 40396 22484 40472 22684
use cut_M1M4_1x2 
transform 1 0 40396 0 1 23444
box 40396 23444 40472 23644
use cut_M1M4_1x2 
transform 1 0 40396 0 1 24404
box 40396 24404 40472 24604
use cut_M1M4_1x2 
transform 1 0 40396 0 1 25364
box 40396 25364 40472 25564
<< labels >>
flabel locali s 40396 0 40696 26808 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 5380 21706 5956 21926 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew
flabel locali s 1060 4058 1636 4278 0 FreeSans 400 0 0 0 VLPF
port 3 nsew
<< end >>
