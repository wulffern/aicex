magic
tech sky130A
magscale 1 2
timestamp 1659354078
<< checkpaint >>
rect 0 0 2520 352
<< locali >>
rect -108 146 540 206
rect 432 146 600 206
rect 600 58 864 118
rect 600 58 660 206
rect 432 146 600 206
rect 600 234 864 294
rect 600 146 660 294
rect 1656 58 1824 118
rect 1824 146 2088 206
rect 1824 58 1884 206
rect 1656 234 1824 294
rect 1824 146 2088 206
rect 1824 146 1884 294
<< m3 >>
rect 756 0 956 352
rect 756 0 956 352
use SUNTRB_NCHDL MN1
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTRB_PCHDL MP1
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 234
box 756 234 956 310
use SUNTRB_cut_M1M4_2x1 
transform 1 0 756 0 1 58
box 756 58 956 134
<< labels >>
flabel m3 s 756 0 956 352 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
<< end >>
