magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 8460 960
<< m1 >>
rect 90 -40 8430 40
rect 8370 40 8430 120
rect 90 120 8310 200
rect 8370 120 8430 200
rect 90 200 150 280
rect 8370 200 8430 280
rect 90 280 150 360
rect 210 280 8430 360
rect 90 360 150 440
rect 8370 360 8430 440
rect 90 440 8310 520
rect 8370 440 8430 520
rect 90 520 150 600
rect 8370 520 8430 600
rect 90 600 150 680
rect 210 600 8430 680
rect 90 680 150 760
rect 90 760 8430 840
<< m2 >>
rect 90 -40 8430 40
rect 8370 40 8430 120
rect 90 120 8310 200
rect 8370 120 8430 200
rect 90 200 150 280
rect 8370 200 8430 280
rect 90 280 150 360
rect 210 280 8430 360
rect 90 360 150 440
rect 8370 360 8430 440
rect 90 440 8310 520
rect 8370 440 8430 520
rect 90 520 150 600
rect 8370 520 8430 600
rect 90 600 150 680
rect 210 600 8430 680
rect 90 680 150 760
rect 90 760 8430 840
<< locali >>
rect 90 -40 8430 40
rect 8370 40 8430 120
rect 90 120 8310 200
rect 8370 120 8430 200
rect 90 200 150 280
rect 8370 200 8430 280
rect 90 280 150 360
rect 210 280 8430 360
rect 90 360 150 440
rect 8370 360 8430 440
rect 90 440 8310 520
rect 8370 440 8430 520
rect 90 520 150 600
rect 8370 520 8430 600
rect 90 600 150 680
rect 210 600 8430 680
rect 90 680 150 760
rect 90 760 8430 840
<< v1 >>
rect 8130 -32 8190 -24
rect 8130 -24 8190 -16
rect 8130 -16 8190 -8
rect 8130 -8 8190 0
rect 8130 0 8190 8
rect 8130 8 8190 16
rect 8130 16 8190 24
rect 8130 24 8190 32
rect 8190 -32 8250 -24
rect 8190 -24 8250 -16
rect 8190 -16 8250 -8
rect 8190 -8 8250 0
rect 8190 0 8250 8
rect 8190 8 8250 16
rect 8190 16 8250 24
rect 8190 24 8250 32
rect 8250 -32 8310 -24
rect 8250 -24 8310 -16
rect 8250 -16 8310 -8
rect 8250 -8 8310 0
rect 8250 0 8310 8
rect 8250 8 8310 16
rect 8250 16 8310 24
rect 8250 24 8310 32
rect 270 128 330 136
rect 270 136 330 144
rect 270 144 330 152
rect 270 152 330 160
rect 270 160 330 168
rect 270 168 330 176
rect 270 176 330 184
rect 270 184 330 192
rect 330 128 390 136
rect 330 136 390 144
rect 330 144 390 152
rect 330 152 390 160
rect 330 160 390 168
rect 330 168 390 176
rect 330 176 390 184
rect 330 184 390 192
rect 390 128 450 136
rect 390 136 450 144
rect 390 144 450 152
rect 390 152 450 160
rect 390 160 450 168
rect 390 168 450 176
rect 390 176 450 184
rect 390 184 450 192
rect 8130 288 8190 296
rect 8130 296 8190 304
rect 8130 304 8190 312
rect 8130 312 8190 320
rect 8130 320 8190 328
rect 8130 328 8190 336
rect 8130 336 8190 344
rect 8130 344 8190 352
rect 8190 288 8250 296
rect 8190 296 8250 304
rect 8190 304 8250 312
rect 8190 312 8250 320
rect 8190 320 8250 328
rect 8190 328 8250 336
rect 8190 336 8250 344
rect 8190 344 8250 352
rect 8250 288 8310 296
rect 8250 296 8310 304
rect 8250 304 8310 312
rect 8250 312 8310 320
rect 8250 320 8310 328
rect 8250 328 8310 336
rect 8250 336 8310 344
rect 8250 344 8310 352
rect 270 448 330 456
rect 270 456 330 464
rect 270 464 330 472
rect 270 472 330 480
rect 270 480 330 488
rect 270 488 330 496
rect 270 496 330 504
rect 270 504 330 512
rect 330 448 390 456
rect 330 456 390 464
rect 330 464 390 472
rect 330 472 390 480
rect 330 480 390 488
rect 330 488 390 496
rect 330 496 390 504
rect 330 504 390 512
rect 390 448 450 456
rect 390 456 450 464
rect 390 464 450 472
rect 390 472 450 480
rect 390 480 450 488
rect 390 488 450 496
rect 390 496 450 504
rect 390 504 450 512
rect 8130 608 8190 616
rect 8130 616 8190 624
rect 8130 624 8190 632
rect 8130 632 8190 640
rect 8130 640 8190 648
rect 8130 648 8190 656
rect 8130 656 8190 664
rect 8130 664 8190 672
rect 8190 608 8250 616
rect 8190 616 8250 624
rect 8190 624 8250 632
rect 8190 632 8250 640
rect 8190 640 8250 648
rect 8190 648 8250 656
rect 8190 656 8250 664
rect 8190 664 8250 672
rect 8250 608 8310 616
rect 8250 616 8310 624
rect 8250 624 8310 632
rect 8250 632 8310 640
rect 8250 640 8310 648
rect 8250 648 8310 656
rect 8250 656 8310 664
rect 8250 664 8310 672
rect 270 768 330 776
rect 270 776 330 784
rect 270 784 330 792
rect 270 792 330 800
rect 270 800 330 808
rect 270 808 330 816
rect 270 816 330 824
rect 270 824 330 832
rect 330 768 390 776
rect 330 776 390 784
rect 330 784 390 792
rect 330 792 390 800
rect 330 800 390 808
rect 330 808 390 816
rect 330 816 390 824
rect 330 824 390 832
rect 390 768 450 776
rect 390 776 450 784
rect 390 784 450 792
rect 390 792 450 800
rect 390 800 450 808
rect 390 808 450 816
rect 390 816 450 824
rect 390 824 450 832
<< v2 >>
rect 8130 -32 8190 -24
rect 8130 -24 8190 -16
rect 8130 -16 8190 -8
rect 8130 -8 8190 0
rect 8130 0 8190 8
rect 8130 8 8190 16
rect 8130 16 8190 24
rect 8130 24 8190 32
rect 8190 -32 8250 -24
rect 8190 -24 8250 -16
rect 8190 -16 8250 -8
rect 8190 -8 8250 0
rect 8190 0 8250 8
rect 8190 8 8250 16
rect 8190 16 8250 24
rect 8190 24 8250 32
rect 8250 -32 8310 -24
rect 8250 -24 8310 -16
rect 8250 -16 8310 -8
rect 8250 -8 8310 0
rect 8250 0 8310 8
rect 8250 8 8310 16
rect 8250 16 8310 24
rect 8250 24 8310 32
rect 270 128 330 136
rect 270 136 330 144
rect 270 144 330 152
rect 270 152 330 160
rect 270 160 330 168
rect 270 168 330 176
rect 270 176 330 184
rect 270 184 330 192
rect 330 128 390 136
rect 330 136 390 144
rect 330 144 390 152
rect 330 152 390 160
rect 330 160 390 168
rect 330 168 390 176
rect 330 176 390 184
rect 330 184 390 192
rect 390 128 450 136
rect 390 136 450 144
rect 390 144 450 152
rect 390 152 450 160
rect 390 160 450 168
rect 390 168 450 176
rect 390 176 450 184
rect 390 184 450 192
rect 8130 288 8190 296
rect 8130 296 8190 304
rect 8130 304 8190 312
rect 8130 312 8190 320
rect 8130 320 8190 328
rect 8130 328 8190 336
rect 8130 336 8190 344
rect 8130 344 8190 352
rect 8190 288 8250 296
rect 8190 296 8250 304
rect 8190 304 8250 312
rect 8190 312 8250 320
rect 8190 320 8250 328
rect 8190 328 8250 336
rect 8190 336 8250 344
rect 8190 344 8250 352
rect 8250 288 8310 296
rect 8250 296 8310 304
rect 8250 304 8310 312
rect 8250 312 8310 320
rect 8250 320 8310 328
rect 8250 328 8310 336
rect 8250 336 8310 344
rect 8250 344 8310 352
rect 270 448 330 456
rect 270 456 330 464
rect 270 464 330 472
rect 270 472 330 480
rect 270 480 330 488
rect 270 488 330 496
rect 270 496 330 504
rect 270 504 330 512
rect 330 448 390 456
rect 330 456 390 464
rect 330 464 390 472
rect 330 472 390 480
rect 330 480 390 488
rect 330 488 390 496
rect 330 496 390 504
rect 330 504 390 512
rect 390 448 450 456
rect 390 456 450 464
rect 390 464 450 472
rect 390 472 450 480
rect 390 480 450 488
rect 390 488 450 496
rect 390 496 450 504
rect 390 504 450 512
rect 8130 608 8190 616
rect 8130 616 8190 624
rect 8130 624 8190 632
rect 8130 632 8190 640
rect 8130 640 8190 648
rect 8130 648 8190 656
rect 8130 656 8190 664
rect 8130 664 8190 672
rect 8190 608 8250 616
rect 8190 616 8250 624
rect 8190 624 8250 632
rect 8190 632 8250 640
rect 8190 640 8250 648
rect 8190 648 8250 656
rect 8190 656 8250 664
rect 8190 664 8250 672
rect 8250 608 8310 616
rect 8250 616 8310 624
rect 8250 624 8310 632
rect 8250 632 8310 640
rect 8250 640 8310 648
rect 8250 648 8310 656
rect 8250 656 8310 664
rect 8250 664 8310 672
rect 270 768 330 776
rect 270 776 330 784
rect 270 784 330 792
rect 270 792 330 800
rect 270 800 330 808
rect 270 808 330 816
rect 270 816 330 824
rect 270 824 330 832
rect 330 768 390 776
rect 330 776 390 784
rect 330 784 390 792
rect 330 792 390 800
rect 330 800 390 808
rect 330 808 390 816
rect 330 816 390 824
rect 330 824 390 832
rect 390 768 450 776
rect 390 776 450 784
rect 390 784 450 792
rect 390 792 450 800
rect 390 800 450 808
rect 390 808 450 816
rect 390 816 450 824
rect 390 824 450 832
<< viali >>
rect 8130 -32 8190 -24
rect 8130 -24 8190 -16
rect 8130 -16 8190 -8
rect 8130 -8 8190 0
rect 8130 0 8190 8
rect 8130 8 8190 16
rect 8130 16 8190 24
rect 8130 24 8190 32
rect 8190 -32 8250 -24
rect 8190 -24 8250 -16
rect 8190 -16 8250 -8
rect 8190 -8 8250 0
rect 8190 0 8250 8
rect 8190 8 8250 16
rect 8190 16 8250 24
rect 8190 24 8250 32
rect 8250 -32 8310 -24
rect 8250 -24 8310 -16
rect 8250 -16 8310 -8
rect 8250 -8 8310 0
rect 8250 0 8310 8
rect 8250 8 8310 16
rect 8250 16 8310 24
rect 8250 24 8310 32
rect 270 128 330 136
rect 270 136 330 144
rect 270 144 330 152
rect 270 152 330 160
rect 270 160 330 168
rect 270 168 330 176
rect 270 176 330 184
rect 270 184 330 192
rect 330 128 390 136
rect 330 136 390 144
rect 330 144 390 152
rect 330 152 390 160
rect 330 160 390 168
rect 330 168 390 176
rect 330 176 390 184
rect 330 184 390 192
rect 390 128 450 136
rect 390 136 450 144
rect 390 144 450 152
rect 390 152 450 160
rect 390 160 450 168
rect 390 168 450 176
rect 390 176 450 184
rect 390 184 450 192
rect 8130 288 8190 296
rect 8130 296 8190 304
rect 8130 304 8190 312
rect 8130 312 8190 320
rect 8130 320 8190 328
rect 8130 328 8190 336
rect 8130 336 8190 344
rect 8130 344 8190 352
rect 8190 288 8250 296
rect 8190 296 8250 304
rect 8190 304 8250 312
rect 8190 312 8250 320
rect 8190 320 8250 328
rect 8190 328 8250 336
rect 8190 336 8250 344
rect 8190 344 8250 352
rect 8250 288 8310 296
rect 8250 296 8310 304
rect 8250 304 8310 312
rect 8250 312 8310 320
rect 8250 320 8310 328
rect 8250 328 8310 336
rect 8250 336 8310 344
rect 8250 344 8310 352
rect 270 448 330 456
rect 270 456 330 464
rect 270 464 330 472
rect 270 472 330 480
rect 270 480 330 488
rect 270 488 330 496
rect 270 496 330 504
rect 270 504 330 512
rect 330 448 390 456
rect 330 456 390 464
rect 330 464 390 472
rect 330 472 390 480
rect 330 480 390 488
rect 330 488 390 496
rect 330 496 390 504
rect 330 504 390 512
rect 390 448 450 456
rect 390 456 450 464
rect 390 464 450 472
rect 390 472 450 480
rect 390 480 450 488
rect 390 488 450 496
rect 390 496 450 504
rect 390 504 450 512
rect 8130 608 8190 616
rect 8130 616 8190 624
rect 8130 624 8190 632
rect 8130 632 8190 640
rect 8130 640 8190 648
rect 8130 648 8190 656
rect 8130 656 8190 664
rect 8130 664 8190 672
rect 8190 608 8250 616
rect 8190 616 8250 624
rect 8190 624 8250 632
rect 8190 632 8250 640
rect 8190 640 8250 648
rect 8190 648 8250 656
rect 8190 656 8250 664
rect 8190 664 8250 672
rect 8250 608 8310 616
rect 8250 616 8310 624
rect 8250 624 8310 632
rect 8250 632 8310 640
rect 8250 640 8310 648
rect 8250 648 8310 656
rect 8250 656 8310 664
rect 8250 664 8310 672
rect 270 768 330 776
rect 270 776 330 784
rect 270 784 330 792
rect 270 792 330 800
rect 270 800 330 808
rect 270 808 330 816
rect 270 816 330 824
rect 270 824 330 832
rect 330 768 390 776
rect 330 776 390 784
rect 330 784 390 792
rect 330 792 390 800
rect 330 800 390 808
rect 330 808 390 816
rect 330 816 390 824
rect 330 824 390 832
rect 390 768 450 776
rect 390 776 450 784
rect 390 784 450 792
rect 390 792 450 800
rect 390 800 450 808
rect 390 808 450 816
rect 390 816 450 824
rect 390 824 450 832
<< m3 >>
rect 90 -40 8430 40
rect 90 -40 8430 40
rect 8370 40 8430 120
rect 90 120 8130 200
rect 8190 120 8310 200
rect 8370 120 8430 200
rect 90 200 150 280
rect 8370 200 8430 280
rect 90 280 150 360
rect 210 280 270 360
rect 330 280 8430 360
rect 90 360 150 440
rect 8370 360 8430 440
rect 90 440 8310 520
rect 8370 440 8430 520
rect 90 520 150 600
rect 8370 520 8430 600
rect 90 600 150 680
rect 210 600 8430 680
rect 90 680 150 760
rect 90 760 8430 840
rect 90 760 8430 840
<< rm3 >>
rect 8130 120 8190 200
rect 270 280 330 360
<< labels >>
flabel m3 s 90 -40 8430 40 0 FreeSans 400 0 0 0 B
port 1 nsew
flabel m3 s 90 760 8430 840 0 FreeSans 400 0 0 0 A
port 2 nsew
<< end >>
