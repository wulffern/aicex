magic
tech sky130A
magscale 1 2
timestamp 1661020682
<< checkpaint >>
rect 0 0 2520 4928
<< locali >>
rect 1656 234 1824 294
rect 1824 790 2040 850
rect 1824 234 1884 850
rect 1980 850 2088 910
rect 1656 938 1824 998
rect 1824 1554 2088 1614
rect 1824 4370 2088 4430
rect 1824 938 1884 4430
rect 432 2258 600 2318
rect 600 938 864 998
rect 600 938 660 2318
rect 480 3254 600 3314
rect 600 938 864 998
rect 600 938 660 3314
rect 432 3314 540 3374
rect 864 1642 1032 1702
rect 864 2346 1032 2406
rect 1032 1642 1092 2406
rect 432 4722 600 4782
rect 600 4458 864 4518
rect 600 4458 660 4782
rect 324 1202 540 1262
rect 324 146 540 206
rect 756 4810 972 4870
rect 756 4458 972 4518
rect 324 3666 540 3726
rect 2412 132 2628 220
rect -108 132 108 220
<< m1 >>
rect 2088 2258 2256 2318
rect 2088 3314 2256 3374
rect 1656 234 2256 294
rect 2256 234 2316 3382
rect 480 1494 600 1554
rect 600 586 864 646
rect 600 586 660 1622
rect 432 1554 540 1614
rect 864 3402 1032 3462
rect 864 4458 1032 4518
rect 1032 3402 1092 4526
rect 432 2610 600 2670
rect 600 2346 864 2406
rect 600 2346 660 2678
rect 1656 2698 1824 2758
rect 1824 1906 2088 1966
rect 1824 2962 2088 3022
rect 1824 1906 1884 3030
rect 1656 4810 1824 4870
rect 1824 4018 2088 4078
rect 1824 4018 1884 4878
rect 204 498 432 558
rect 204 3666 432 3726
rect 204 498 264 3734
<< m2 >>
rect 432 4370 604 4446
rect 604 3314 2088 3390
rect 604 3314 680 4446
<< m3 >>
rect 1548 0 1748 4928
rect 756 0 956 4928
rect 1548 0 1748 4928
rect 756 0 956 4928
use SUNTRB_ XA0
transform 1 0 0 0 1 0
box 0 0 0 0
use SUNTRB_NDX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2520 704
use SUNTRB_IVX1_CV XA2
transform 1 0 0 0 1 704
box 0 704 2520 1056
use SUNTRB_IVTRIX1_CV XA3
transform 1 0 0 0 1 1056
box 0 1056 2520 1760
use SUNTRB_IVTRIX1_CV XA4
transform 1 0 0 0 1 1760
box 0 1760 2520 2464
use SUNTRB_IVX1_CV XA5
transform 1 0 0 0 1 2464
box 0 2464 2520 2816
use SUNTRB_IVTRIX1_CV XA6
transform 1 0 0 0 1 2816
box 0 2816 2520 3520
use SUNTRB_NDTRIX1_CV XA7
transform 1 0 0 0 1 3520
box 0 3520 2520 4576
use SUNTRB_IVX1_CV XA8
transform 1 0 0 0 1 4576
box 0 4576 2520 4928
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1980 0 1 2258
box 1980 2258 2164 2326
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1980 0 1 3314
box 1980 3314 2164 3382
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1548 0 1 234
box 1548 234 1732 302
use SUNTRB_cut_M1M2_2x1 
transform 1 0 324 0 1 1554
box 324 1554 508 1622
use SUNTRB_cut_M1M2_2x1 
transform 1 0 756 0 1 586
box 756 586 940 654
use SUNTRB_cut_M1M3_2x1 
transform 1 0 324 0 1 4370
box 324 4370 524 4446
use SUNTRB_cut_M1M3_2x1 
transform 1 0 1980 0 1 3314
box 1980 3314 2180 3390
use SUNTRB_cut_M1M2_2x1 
transform 1 0 756 0 1 3402
box 756 3402 940 3470
use SUNTRB_cut_M1M2_2x1 
transform 1 0 756 0 1 4458
box 756 4458 940 4526
use SUNTRB_cut_M1M2_2x1 
transform 1 0 324 0 1 2610
box 324 2610 508 2678
use SUNTRB_cut_M1M2_2x1 
transform 1 0 756 0 1 2346
box 756 2346 940 2414
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1548 0 1 2698
box 1548 2698 1732 2766
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1980 0 1 1906
box 1980 1906 2164 1974
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1980 0 1 2962
box 1980 2962 2164 3030
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1548 0 1 4810
box 1548 4810 1732 4878
use SUNTRB_cut_M1M2_2x1 
transform 1 0 1980 0 1 4018
box 1980 4018 2164 4086
use SUNTRB_cut_M1M2_2x1 
transform 1 0 324 0 1 498
box 324 498 508 566
use SUNTRB_cut_M1M2_2x1 
transform 1 0 324 0 1 3666
box 324 3666 508 3734
<< labels >>
flabel locali s 324 1202 540 1262 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 CK
port 2 nsew
flabel locali s 756 4810 972 4870 0 FreeSans 400 0 0 0 Q
port 4 nsew
flabel locali s 756 4458 972 4518 0 FreeSans 400 0 0 0 QN
port 5 nsew
flabel locali s 324 3666 540 3726 0 FreeSans 400 0 0 0 RN
port 3 nsew
flabel locali s 2412 132 2628 220 0 FreeSans 400 0 0 0 BULKP
port 6 nsew
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 BULKN
port 7 nsew
flabel m3 s 1548 0 1748 4928 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 756 0 956 4928 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
