magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 13120
<< locali >>
rect 360 5250 514 5310
rect 514 4050 720 4110
rect 514 4050 574 5310
rect 360 7810 514 7870
rect 514 6610 720 6670
rect 514 6610 574 7870
rect 1526 3970 1740 4030
rect 1380 3730 1526 3790
rect 1526 3730 1586 4030
rect 360 10690 514 10750
rect 514 10450 720 10510
rect 514 10450 574 10750
rect 330 10690 390 11070
rect 390 11590 514 11650
rect 514 11410 720 11470
rect 514 11410 574 11650
rect 390 11650 450 11710
rect 390 11910 514 11970
rect 514 11730 720 11790
rect 514 11730 574 11970
rect 390 11970 450 12030
rect 360 12610 514 12670
rect 514 12210 720 12270
rect 514 12210 574 12670
rect 1380 7890 1534 7950
rect 1534 9090 1740 9150
rect 1534 7890 1594 9150
rect 1650 3650 1830 3710
rect 270 3010 450 3070
rect 270 12290 450 12350
rect 1290 12690 1470 12750
rect 270 9410 450 9470
rect 630 10770 810 10830
<< m1 >>
rect 360 6530 514 6590
rect 514 2770 720 2830
rect 514 2770 574 6598
rect 1740 10370 1894 10430
rect 1380 690 1894 750
rect 1894 690 1954 10438
rect 360 11330 514 11390
rect 514 10130 720 10190
rect 514 10130 574 11398
rect 1380 5330 1534 5390
rect 1534 9730 1740 9790
rect 1534 5330 1594 9798
<< m3 >>
rect 1828 4370 1896 8394
rect 266 5246 450 5314
rect 878 5268 946 5452
rect 1014 6548 1082 6732
rect 1150 7828 1218 8012
rect 1770 4370 1954 4554
rect 1290 0 1474 13120
rect 630 0 814 13120
rect 1290 0 1474 13120
rect 630 0 814 13120
<< m2 >>
rect 266 2046 450 2114
rect 266 446 450 514
rect 1286 686 1470 754
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use SARMRYX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2100 3840
use SWX4_CV XA2
transform 1 0 0 0 1 3840
box 0 3840 2100 5120
use SWX4_CV XA3
transform 1 0 0 0 1 5120
box 0 5120 2100 6400
use SWX4_CV XA4
transform 1 0 0 0 1 6400
box 0 6400 2100 7680
use SWX4_CV XA5
transform 1 0 0 0 1 7680
box 0 7680 2100 8960
use SARCEX1_CV XA6
transform 1 0 0 0 1 8960
box 0 8960 2100 10240
use IVX1_CV XA7
transform 1 0 0 0 1 10240
box 0 10240 2100 10560
use IVX1_CV XA8
transform 1 0 0 0 1 10560
box 0 10560 2100 10880
use NDX1_CV XA9
transform 1 0 0 0 1 10880
box 0 10880 2100 11520
use IVX1_CV XA10
transform 1 0 0 0 1 11520
box 0 11520 2100 11840
use NRX1_CV XA11
transform 1 0 0 0 1 11840
box 0 11840 2100 12480
use IVX1_CV XA12
transform 1 0 0 0 1 12480
box 0 12480 2100 12800
use TAPCELLB_CV XA13
transform 1 0 0 0 1 12800
box 0 12800 2100 13120
use DMY_CV XA14
transform 1 0 0 0 1 13120
box 0 13120 0 13120
use cut_M1M2_2x1 
transform 1 0 270 0 1 6530
box 270 6530 454 6598
use cut_M1M2_2x1 
transform 1 0 630 0 1 2770
box 630 2770 814 2838
use cut_M1M2_2x1 
transform 1 0 1650 0 1 10370
box 1650 10370 1834 10438
use cut_M1M2_2x1 
transform 1 0 1290 0 1 690
box 1290 690 1474 758
use cut_M1M2_2x1 
transform 1 0 270 0 1 11330
box 270 11330 454 11398
use cut_M1M2_2x1 
transform 1 0 630 0 1 10130
box 630 10130 814 10198
use cut_M1M2_2x1 
transform 1 0 1290 0 1 5330
box 1290 5330 1474 5398
use cut_M1M2_2x1 
transform 1 0 1650 0 1 9730
box 1650 9730 1834 9798
use cut_M1M4_2x1 
transform 1 0 266 0 1 5246
box 266 5246 450 5314
use cut_M1M4_1x2 
transform 1 0 878 0 1 5268
box 878 5268 946 5452
use cut_M1M4_1x2 
transform 1 0 1014 0 1 6548
box 1014 6548 1082 6732
use cut_M1M4_1x2 
transform 1 0 1150 0 1 7828
box 1150 7828 1218 8012
use cut_M2M3_2x1 
transform 1 0 1286 0 1 686
box 1286 686 1470 754
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
<< labels >>
flabel m2 s 266 2046 450 2114 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1650 3650 1830 3710 0 FreeSans 400 0 0 0 RST_N
port 2 nsew
flabel m2 s 266 446 450 514 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 270 3010 450 3070 0 FreeSans 400 0 0 0 CMP_ON
port 4 nsew
flabel m2 s 1286 686 1470 754 0 FreeSans 400 0 0 0 ENO
port 5 nsew
flabel m3 s 266 5246 450 5314 0 FreeSans 400 0 0 0 CN1
port 6 nsew
flabel m3 s 878 5268 946 5452 0 FreeSans 400 0 0 0 CP1
port 7 nsew
flabel m3 s 1014 6548 1082 6732 0 FreeSans 400 0 0 0 CP0
port 8 nsew
flabel m3 s 1150 7828 1218 8012 0 FreeSans 400 0 0 0 CN0
port 9 nsew
flabel locali s 270 12290 450 12350 0 FreeSans 400 0 0 0 CEIN
port 10 nsew
flabel locali s 1290 12690 1470 12750 0 FreeSans 400 0 0 0 CEO
port 11 nsew
flabel locali s 270 9410 450 9470 0 FreeSans 400 0 0 0 CKS
port 12 nsew
flabel locali s 630 10770 810 10830 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 1770 4370 1954 4554 0 FreeSans 400 0 0 0 VREF
port 14 nsew
flabel m3 s 1290 0 1474 13120 0 FreeSans 400 0 0 0 AVDD
port 15 nsew
flabel m3 s 630 0 814 13120 0 FreeSans 400 0 0 0 AVSS
port 16 nsew
<< end >>
