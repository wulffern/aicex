magic
tech sky130A
magscale 1 2
timestamp 1661001370
<< checkpaint >>
rect -1560 -1920 47020 41968
<< locali >>
rect 46252 -1392 46492 41440
rect -1032 -1392 46492 -1152
rect -1032 41200 46492 41440
rect -1032 -1392 -792 41440
rect 46252 -1392 46492 41440
rect 46780 -1920 47020 41968
rect -1560 -1920 47020 -1680
rect -1560 41728 47020 41968
rect -1560 -1920 -1320 41968
rect 46780 -1920 47020 41968
rect 15376 6192 29512 6252
rect 38980 26626 39196 26686
rect 26548 498 26764 558
rect 684 146 900 206
use SUN_PLL_BUF xb1
transform 1 0 360 0 1 0
box 360 0 15072 11040
use SUN_PLL_LPF xb2
transform 1 0 360 0 1 11920
box 360 11920 39904 40048
use SUN_PLL_DIVN xc1
transform 1 0 16144 0 1 0
box 16144 0 30280 7020
use SUN_PLL_ROSC xd1
transform 1 0 30640 0 1 0
box 30640 0 37216 5408
use SUN_PLL_KICK xk1
transform 1 0 38656 0 1 0
box 38656 0 42712 14208
use SUN_PLL_CP xk2
transform 1 0 38656 0 1 15088
box 38656 15088 43072 25776
use SUN_PLL_PFD xk3
transform 1 0 38656 0 1 25776
box 38656 25776 42712 31536
use SUN_PLL_BIAS xl1
transform 1 0 43072 0 1 0
box 43072 0 45100 18720
<< labels >>
flabel locali s 46252 -1392 46492 41440 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 46780 -1920 47020 41968 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 15376 6192 29512 6252 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel locali s 38980 26626 39196 26686 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel locali s 26548 498 26764 558 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel locali s 684 146 900 206 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
