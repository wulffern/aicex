magic
tech sky130A
magscale 1 2
timestamp 1658699483
<< checkpaint >>
rect -2284 0 26372 50262
<< m3 >>
rect 9100 28760 26178 28836
rect 9100 29148 26178 29224
rect 24104 29528 24180 37032
rect 24384 29528 24460 44776
rect 3944 29612 4020 40544
rect 4824 29806 4900 40544
rect 8984 30000 9060 40544
rect -216 30194 -140 40544
rect -216 30194 -140 40544
rect 13432 30388 13508 40570
rect 13432 30388 13508 40570
rect 18472 30582 18548 40570
rect 18472 30582 18548 40570
rect 10579 30776 10655 40570
rect 10579 30776 10655 40570
rect 15619 30970 15695 40570
rect 15619 30970 15695 40570
rect 499 31164 575 40570
rect 5539 31358 5615 40570
rect 5539 31358 5615 40570
rect 3352 31552 3428 40570
rect 3352 31552 3428 40570
rect 8392 31746 8468 40570
rect 8392 31746 8468 40570
rect 659 31940 735 41978
rect 8232 32134 8308 41978
rect 5699 32328 5775 41978
rect 3192 32522 3268 41978
rect 10914 32716 10990 43386
rect 13098 32910 13174 43386
rect 15954 33104 16030 43386
rect 8058 33298 8134 43386
rect 3018 33492 3094 43386
rect 834 33686 910 43386
rect 18138 33880 18214 43386
rect 5874 34074 5950 43386
rect 11072 50 11272 126
rect 12816 50 13016 126
rect 20659 40570 20735 40770
rect 1568 39584 1768 39784
rect 8856 0 9056 5280
rect 9648 0 9848 5280
<< m2 >>
rect 14872 28254 14948 28836
rect 9100 28254 9176 29224
rect 3944 29536 14020 29612
rect 4824 29730 13660 29806
rect 8984 29924 13300 30000
rect -216 30118 14380 30194
rect 11304 30312 13508 30388
rect 11664 30506 18548 30582
rect 10579 30700 11200 30776
rect 11484 30894 15695 30970
rect 499 31088 9760 31164
rect 5539 31282 10480 31358
rect 3352 31476 10120 31552
rect 8392 31670 10840 31746
rect 659 31864 9940 31940
rect 8232 32058 11020 32134
rect 5699 32252 10660 32328
rect 3192 32446 10300 32522
rect 10914 32640 12940 32716
rect 12684 32834 13174 32910
rect 12504 33028 16030 33104
rect 8058 33222 13120 33298
rect 3018 33416 13840 33492
rect 834 33610 14200 33686
rect 12324 33804 18214 33880
rect 5874 33998 13480 34074
rect -216 35264 -16 35340
<< m4 >>
rect 24104 29148 24180 29528
rect 24384 28760 24460 29528
<< m1 >>
rect 13944 28194 14020 29536
rect 13584 28194 13660 29730
rect 13224 28194 13300 29924
rect 14304 28194 14380 30118
rect 11304 28194 11380 30312
rect 11664 28194 11740 30506
rect 11124 28194 11200 30700
rect 11484 28194 11560 30894
rect 9684 28194 9760 31088
rect 10404 28194 10480 31282
rect 10044 28194 10120 31476
rect 10764 28194 10840 31670
rect 9864 28194 9940 31864
rect 10944 28194 11020 32058
rect 10584 28194 10660 32252
rect 10224 28194 10300 32446
rect 12864 28194 12940 32640
rect 12684 28194 12760 32834
rect 12504 28194 12580 33028
rect 13044 28194 13120 33222
rect 13764 28194 13840 33416
rect 14124 28194 14200 33610
rect 12324 28194 12400 33804
rect 13404 28194 13480 33998
<< locali >>
rect 11072 2698 11288 2758
rect 11072 1290 11288 1350
rect 20360 46624 20576 46684
rect -232 45128 -16 45188
rect 10064 498 10280 558
use SARBSSW_CV XB1
transform -1 0 12044 0 1 0
box 12044 0 26372 5280
use SARBSSW_CV XB2
transform 1 0 12044 0 1 0
box 12044 0 26372 5280
use CDAC8_CV XDAC1
transform -1 0 11844 0 1 5474
box 11844 5474 23576 28254
use CDAC8_CV XDAC2
transform 1 0 12204 0 1 5474
box 12204 5474 23936 28254
use SARDIGEX4_CV XA0
transform 1 0 -556 0 1 34774
box -556 34774 1964 49206
use SARDIGEX4_CV XA1
transform -1 0 4484 0 1 34774
box 4484 34774 7004 49206
use SARDIGEX4_CV XA2
transform 1 0 4484 0 1 34774
box 4484 34774 7004 49206
use SARDIGEX4_CV XA3
transform -1 0 9524 0 1 34774
box 9524 34774 12044 49206
use SARDIGEX4_CV XA4
transform 1 0 9524 0 1 34774
box 9524 34774 12044 49206
use SARDIGEX4_CV XA5
transform -1 0 14564 0 1 34774
box 14564 34774 17084 49206
use SARDIGEX4_CV XA6
transform 1 0 14564 0 1 34774
box 14564 34774 17084 49206
use SARDIGEX4_CV XA7
transform -1 0 19604 0 1 34774
box 19604 34774 22124 49206
use SARDIGEX4_CV XA8
transform 1 0 19604 0 1 34774
box 19604 34774 22124 49206
use SARCMPX1_CV XA20
transform -1 0 24644 0 1 34774
box 24644 34774 27164 50262
use cut_M3M4_1x2 
transform 1 0 14872 0 1 28254
box 14872 28254 14948 28454
use cut_M3M4_2x1 
transform 1 0 14872 0 1 28760
box 14872 28760 15072 28836
use cut_M3M4_1x2 
transform 1 0 9100 0 1 28254
box 9100 28254 9176 28454
use cut_M3M4_2x1 
transform 1 0 9100 0 1 29148
box 9100 29148 9300 29224
use cut_M2M4_2x1 
transform 1 0 24104 0 1 37032
box 24104 37032 24304 37108
use cut_M4M5_2x1 
transform 1 0 24104 0 1 29148
box 24104 29148 24304 29224
use cut_M4M5_1x2 
transform 1 0 24104 0 1 29528
box 24104 29528 24180 29728
use cut_M3M4_2x1 
transform 1 0 24260 0 1 44776
box 24260 44776 24460 44852
use cut_M2M3_2x1 
transform 1 0 24104 0 1 44776
box 24104 44776 24304 44852
use cut_M4M5_2x1 
transform 1 0 24384 0 1 28760
box 24384 28760 24584 28836
use cut_M4M5_1x2 
transform 1 0 24384 0 1 29528
box 24384 29528 24460 29728
use cut_M3M4_1x2 
transform 1 0 3944 0 1 29474
box 3944 29474 4020 29674
use cut_M2M3_1x2 
transform 1 0 13936 0 1 29474
box 13936 29474 14012 29674
use cut_M3M4_1x2 
transform 1 0 4824 0 1 29668
box 4824 29668 4900 29868
use cut_M2M3_1x2 
transform 1 0 13576 0 1 29668
box 13576 29668 13652 29868
use cut_M3M4_1x2 
transform 1 0 8984 0 1 29862
box 8984 29862 9060 30062
use cut_M2M3_1x2 
transform 1 0 13216 0 1 29862
box 13216 29862 13292 30062
use cut_M3M4_1x2 
transform 1 0 -216 0 1 30056
box -216 30056 -140 30256
use cut_M2M3_1x2 
transform 1 0 14296 0 1 30056
box 14296 30056 14372 30256
use cut_M3M4_1x2 
transform 1 0 13432 0 1 30250
box 13432 30250 13508 30450
use cut_M2M3_1x2 
transform 1 0 11296 0 1 30250
box 11296 30250 11372 30450
use cut_M3M4_1x2 
transform 1 0 18472 0 1 30444
box 18472 30444 18548 30644
use cut_M2M3_1x2 
transform 1 0 11656 0 1 30444
box 11656 30444 11732 30644
use cut_M3M4_1x2 
transform 1 0 10579 0 1 30638
box 10579 30638 10655 30838
use cut_M2M3_1x2 
transform 1 0 11116 0 1 30638
box 11116 30638 11192 30838
use cut_M3M4_1x2 
transform 1 0 15619 0 1 30832
box 15619 30832 15695 31032
use cut_M2M3_1x2 
transform 1 0 11476 0 1 30832
box 11476 30832 11552 31032
use cut_M3M4_1x2 
transform 1 0 499 0 1 31026
box 499 31026 575 31226
use cut_M2M3_1x2 
transform 1 0 9676 0 1 31026
box 9676 31026 9752 31226
use cut_M3M4_1x2 
transform 1 0 5539 0 1 31220
box 5539 31220 5615 31420
use cut_M2M3_1x2 
transform 1 0 10396 0 1 31220
box 10396 31220 10472 31420
use cut_M3M4_1x2 
transform 1 0 3352 0 1 31414
box 3352 31414 3428 31614
use cut_M2M3_1x2 
transform 1 0 10036 0 1 31414
box 10036 31414 10112 31614
use cut_M3M4_1x2 
transform 1 0 8392 0 1 31608
box 8392 31608 8468 31808
use cut_M2M3_1x2 
transform 1 0 10756 0 1 31608
box 10756 31608 10832 31808
use cut_M3M4_1x2 
transform 1 0 659 0 1 31802
box 659 31802 735 32002
use cut_M2M3_1x2 
transform 1 0 9856 0 1 31802
box 9856 31802 9932 32002
use cut_M3M4_1x2 
transform 1 0 8232 0 1 31996
box 8232 31996 8308 32196
use cut_M2M3_1x2 
transform 1 0 10936 0 1 31996
box 10936 31996 11012 32196
use cut_M3M4_1x2 
transform 1 0 5699 0 1 32190
box 5699 32190 5775 32390
use cut_M2M3_1x2 
transform 1 0 10576 0 1 32190
box 10576 32190 10652 32390
use cut_M3M4_1x2 
transform 1 0 3192 0 1 32384
box 3192 32384 3268 32584
use cut_M2M3_1x2 
transform 1 0 10216 0 1 32384
box 10216 32384 10292 32584
use cut_M3M4_1x2 
transform 1 0 10914 0 1 32578
box 10914 32578 10990 32778
use cut_M2M3_1x2 
transform 1 0 12856 0 1 32578
box 12856 32578 12932 32778
use cut_M3M4_1x2 
transform 1 0 13098 0 1 32772
box 13098 32772 13174 32972
use cut_M2M3_1x2 
transform 1 0 12676 0 1 32772
box 12676 32772 12752 32972
use cut_M3M4_1x2 
transform 1 0 15954 0 1 32966
box 15954 32966 16030 33166
use cut_M2M3_1x2 
transform 1 0 12496 0 1 32966
box 12496 32966 12572 33166
use cut_M3M4_1x2 
transform 1 0 8058 0 1 33160
box 8058 33160 8134 33360
use cut_M2M3_1x2 
transform 1 0 13036 0 1 33160
box 13036 33160 13112 33360
use cut_M3M4_1x2 
transform 1 0 3018 0 1 33354
box 3018 33354 3094 33554
use cut_M2M3_1x2 
transform 1 0 13756 0 1 33354
box 13756 33354 13832 33554
use cut_M3M4_1x2 
transform 1 0 834 0 1 33548
box 834 33548 910 33748
use cut_M2M3_1x2 
transform 1 0 14116 0 1 33548
box 14116 33548 14192 33748
use cut_M3M4_1x2 
transform 1 0 18138 0 1 33742
box 18138 33742 18214 33942
use cut_M2M3_1x2 
transform 1 0 12316 0 1 33742
box 12316 33742 12392 33942
use cut_M3M4_1x2 
transform 1 0 5874 0 1 33936
box 5874 33936 5950 34136
use cut_M2M3_1x2 
transform 1 0 13396 0 1 33936
box 13396 33936 13472 34136
<< labels >>
flabel m3 s -216 30194 -140 40544 0 FreeSans 400 0 0 0 D<8>
port 6 nsew
flabel m3 s 13432 30388 13508 40570 0 FreeSans 400 0 0 0 D<3>
port 11 nsew
flabel m3 s 18472 30582 18548 40570 0 FreeSans 400 0 0 0 D<1>
port 13 nsew
flabel m3 s 10579 30776 10655 40570 0 FreeSans 400 0 0 0 D<4>
port 10 nsew
flabel m3 s 15619 30970 15695 40570 0 FreeSans 400 0 0 0 D<2>
port 12 nsew
flabel m3 s 5539 31358 5615 40570 0 FreeSans 400 0 0 0 D<6>
port 8 nsew
flabel m3 s 3352 31552 3428 40570 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8392 31746 8468 40570 0 FreeSans 400 0 0 0 D<5>
port 9 nsew
flabel m3 s 11072 50 11272 126 0 FreeSans 400 0 0 0 SAR_IP
port 1 nsew
flabel m3 s 12816 50 13016 126 0 FreeSans 400 0 0 0 SAR_IN
port 2 nsew
flabel locali s 11072 2698 11288 2758 0 FreeSans 400 0 0 0 SARN
port 3 nsew
flabel locali s 11072 1290 11288 1350 0 FreeSans 400 0 0 0 SARP
port 4 nsew
flabel locali s 20360 46624 20576 46684 0 FreeSans 400 0 0 0 DONE
port 5 nsew
flabel m3 s 20659 40570 20735 40770 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
flabel m2 s -216 35264 -16 35340 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s -232 45128 -16 45188 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 10064 498 10280 558 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel m3 s 1568 39584 1768 39784 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel m3 s 8856 0 9056 5280 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel m3 s 9648 0 9848 5280 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
<< end >>
