magic
tech sky130A
magscale 1 2
timestamp 1660085871
<< checkpaint >>
rect 0 -896 43334 14320
<< m2 >>
rect 11902 -896 25078 -592
rect 0 -592 11520 -288
<< locali >>
rect 25694 -204 43334 -144
rect 31526 7890 31742 7950
rect 41138 498 41354 558
rect 12226 146 12442 206
use SUN_PLL_LPF xa1
transform 1 0 0 0 1 0
box 0 0 11614 14320
use SUN_PLL_BUF xb1
transform 1 0 11902 0 1 0
box 11902 0 25406 11456
use SUN_PLL_DIVN xh1
transform 1 0 25694 0 1 0
box 25694 0 43334 6958
use SUN_PLL_ROSC xh2
transform 1 0 25694 0 1 6958
box 25694 6958 30842 11550
use SUN_PLL_PFD xj1
transform 1 0 31202 0 1 7040
box 31202 7040 33722 10912
use SUN_PLL_CP xk1
transform 1 0 34010 0 1 7040
box 34010 7040 36530 11808
use SUN_PLL_BIAS xl2
transform 1 0 36818 0 1 7040
box 36818 7040 39446 10928
<< labels >>
flabel m2 s 11902 -896 25078 -592 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 0 -592 11520 -288 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 25694 -204 43334 -144 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel locali s 31526 7890 31742 7950 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel locali s 41138 498 41354 558 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel locali s 12226 146 12442 206 0 FreeSans 400 0 0 0 IBSPR_1U
port 6 nsew
<< end >>
