magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 4416 7696
<< locali >>
rect 3792 384 4032 7312
rect 384 384 4032 624
rect 384 7072 4032 7312
rect 384 384 624 7312
rect 3792 384 4032 7312
rect 4176 0 4416 7696
rect 0 0 4416 240
rect 0 7456 4416 7696
rect 0 0 240 7696
rect 4176 0 4416 7696
rect 1632 2410 1800 2470
rect 1632 2586 1800 2646
rect 1632 3114 1800 3174
rect 1800 2410 1860 3174
rect 3252 826 3420 886
rect 3252 2058 3420 2118
rect 3252 3290 3420 3350
rect 3252 4522 3420 4582
rect 3252 5754 3420 5814
rect 3420 826 3480 5814
<< m1 >>
rect 1524 384 1740 886
rect 660 384 876 988
rect 660 384 876 2748
rect 660 384 876 3276
rect 3144 0 3360 886
rect 2280 0 2496 988
rect 2820 5842 2988 5902
rect 2988 1002 3252 1062
rect 2820 3378 2988 3438
rect 2820 4610 2988 4670
rect 1632 3290 2988 3350
rect 2988 1002 3048 5902
<< m2 >>
rect 2820 914 2992 990
rect 1632 2762 2992 2838
rect 2992 2234 3252 2310
rect 2820 2146 2992 2222
rect 2992 914 3068 2838
rect 0 2674 216 2734
rect 0 3202 216 3262
rect 0 3466 216 3526
rect 0 914 216 974
rect 0 914 216 974
rect 952 914 1200 990
rect 108 914 952 990
rect 952 914 1028 990
rect 0 2674 216 2734
rect 952 2674 1200 2750
rect 108 2674 952 2750
rect 952 2674 1028 2750
rect 0 3202 216 3262
rect 952 3202 1200 3278
rect 108 3202 952 3278
rect 952 3202 1028 3278
rect 0 3466 216 3526
rect 3004 3466 3252 3542
rect 108 3466 3004 3542
rect 3004 3466 3080 3542
<< m3 >>
rect 3252 3466 3432 3542
rect 3252 4698 3432 4774
rect 3252 5930 3432 6006
rect 3432 3466 3508 6006
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa10
transform 1 0 768 0 1 768
box 768 768 2028 2528
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa20
transform 1 0 768 0 1 2528
box 768 2528 2028 3056
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa40
transform 1 0 768 0 1 3056
box 768 3056 2028 3584
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc10
transform -1 0 3648 0 1 768
box 3648 768 4908 2000
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc20
transform -1 0 3648 0 1 2000
box 3648 2000 4908 3232
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_00
transform -1 0 3648 0 1 3232
box 3648 3232 4908 4464
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_10
transform -1 0 3648 0 1 4464
box 3648 4464 4908 5696
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_20
transform -1 0 3648 0 1 5696
box 3648 5696 4908 6928
use cut_M1M2_2x1 
transform 1 0 1540 0 1 826
box 1540 826 1724 894
use cut_M1M2_2x1 
transform 1 0 1540 0 1 384
box 1540 384 1724 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 900
box 676 900 860 968
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 2660
box 676 2660 860 2728
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 3188
box 676 3188 860 3256
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 3160 0 1 826
box 3160 826 3344 894
use cut_M1M2_2x1 
transform 1 0 3160 0 1 0
box 3160 0 3344 68
use cut_M1M2_2x1 
transform 1 0 2296 0 1 900
box 2296 900 2480 968
use cut_M1M2_2x1 
transform 1 0 2296 0 1 0
box 2296 0 2480 68
use cut_M1M2_2x1 
transform 1 0 2712 0 1 5842
box 2712 5842 2896 5910
use cut_M1M2_2x1 
transform 1 0 3144 0 1 1002
box 3144 1002 3328 1070
use cut_M1M2_2x1 
transform 1 0 2712 0 1 3378
box 2712 3378 2896 3446
use cut_M1M2_2x1 
transform 1 0 2712 0 1 4610
box 2712 4610 2896 4678
use cut_M1M2_2x1 
transform 1 0 1524 0 1 3290
box 1524 3290 1708 3358
use cut_M1M3_2x1 
transform 1 0 2712 0 1 914
box 2712 914 2912 990
use cut_M1M3_2x1 
transform 1 0 1524 0 1 2762
box 1524 2762 1724 2838
use cut_M1M3_2x1 
transform 1 0 3144 0 1 2234
box 3144 2234 3344 2310
use cut_M1M3_2x1 
transform 1 0 2712 0 1 2146
box 2712 2146 2912 2222
use cut_M1M4_2x1 
transform 1 0 3144 0 1 3466
box 3144 3466 3344 3542
use cut_M1M4_2x1 
transform 1 0 3144 0 1 4698
box 3144 4698 3344 4774
use cut_M1M4_2x1 
transform 1 0 3144 0 1 5930
box 3144 5930 3344 6006
use cut_M1M3_2x1 
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M3_2x1 
transform 1 0 1108 0 1 2674
box 1108 2674 1308 2750
use cut_M1M3_2x1 
transform 1 0 1108 0 1 3202
box 1108 3202 1308 3278
use cut_M1M3_2x1 
transform 1 0 3160 0 1 3466
box 3160 3466 3360 3542
<< labels >>
flabel locali s 3792 384 4032 7312 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 4176 0 4416 7696 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 0 2674 216 2734 0 FreeSans 400 0 0 0 VFB
port 2 nsew
flabel m2 s 0 3202 216 3262 0 FreeSans 400 0 0 0 VI
port 3 nsew
flabel m2 s 0 3466 216 3526 0 FreeSans 400 0 0 0 VO
port 4 nsew
flabel m2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew
<< end >>
