magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 1050 320
<< pdiff >>
rect 240 40 420 120
rect 240 120 420 200
rect 240 200 420 280
<< ntap >>
rect 960 -40 1140 40
rect 960 40 1140 120
rect 960 120 1140 200
rect 960 200 1140 280
rect 960 280 1140 360
<< poly >>
rect 180 -18 780 18
rect 180 142 780 178
rect 180 302 780 338
rect 600 120 780 200
<< locali >>
rect 600 130 780 190
rect 960 -40 1140 40
rect 240 50 420 110
rect 240 50 420 110
rect 960 40 1140 120
rect 600 130 780 190
rect 960 120 1140 200
rect 960 120 1140 200
rect 240 210 420 270
rect 240 210 420 270
rect 960 200 1140 280
rect 960 280 1140 360
<< pcontact >>
rect 620 140 660 160
rect 620 160 660 180
rect 660 140 720 160
rect 660 160 720 180
rect 720 140 760 160
rect 720 160 760 180
<< ntapc >>
rect 1020 40 1080 120
rect 1020 120 1080 200
rect 1020 200 1080 280
<< pdcontact >>
rect 260 60 300 80
rect 260 80 300 100
rect 300 60 360 80
rect 300 80 360 100
rect 360 60 400 80
rect 360 80 400 100
rect 260 220 300 240
rect 260 240 300 260
rect 300 220 360 240
rect 300 240 360 260
rect 360 220 400 240
rect 360 240 400 260
<< nwell >>
rect 0 -120 1200 440
<< labels >>
flabel locali s 600 130 780 190 0 FreeSans 400 0 0 0 G
port 1 nsew
flabel locali s 240 50 420 110 0 FreeSans 400 0 0 0 S
port 2 nsew
flabel locali s 960 120 1140 200 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 240 210 420 270 0 FreeSans 400 0 0 0 D
port 4 nsew
<< end >>
