magic
tech sky130A
magscale 1 2
timestamp 1660036205
<< checkpaint >>
rect 0 0 200 76
<< m1 >>
rect 0 0 184 68
<< m2 >>
rect 0 0 200 76
<< v1 >>
rect 12 6 172 62
<< labels >>
<< end >>
