magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 960
<< locali >>
rect 720 50 874 110
rect 874 50 1380 110
rect 874 50 934 110
rect 720 850 874 910
rect 874 850 1380 910
rect 874 850 934 910
rect 720 690 874 750
rect 874 690 1380 750
rect 874 690 934 750
rect 330 130 390 510
rect 360 770 514 830
rect 514 50 720 110
rect 514 50 574 830
rect 1740 130 1894 190
rect 1740 770 1894 830
rect 1894 130 1954 830
rect 690 210 750 430
rect 690 530 750 750
rect 1350 210 1410 430
rect 1350 530 1410 750
rect 1650 130 1830 190
rect 1290 690 1470 750
rect 630 850 810 910
<< poly >>
rect 270 142 1830 178
<< m3 >>
rect 1380 370 1534 438
rect 1534 450 1740 518
rect 1534 370 1602 518
rect 1290 0 1474 960
rect 630 0 814 960
rect 1290 0 1474 960
rect 630 0 814 960
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1050 960
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1_DMY
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL MP2
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use cut_M1M4_2x1 
transform 1 0 1290 0 1 370
box 1290 370 1474 438
use cut_M1M4_2x1 
transform 1 0 1650 0 1 450
box 1650 450 1834 518
use cut_M1M4_2x1 
transform 1 0 1290 0 1 210
box 1290 210 1474 278
use cut_M1M4_2x1 
transform 1 0 630 0 1 210
box 630 210 814 278
use cut_M1M4_2x1 
transform 1 0 630 0 1 370
box 630 370 814 438
<< labels >>
flabel locali s 1650 130 1830 190 0 FreeSans 400 0 0 0 C
port 1 nsew
flabel locali s 1290 690 1470 750 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 630 850 810 910 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel m3 s 1290 0 1474 960 0 FreeSans 400 0 0 0 AVDD
port 4 nsew
flabel m3 s 630 0 814 960 0 FreeSans 400 0 0 0 AVSS
port 5 nsew
<< end >>
