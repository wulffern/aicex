magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 1280
<< locali >>
rect 800 1170 968 1230
rect 968 50 1520 110
rect 968 1170 1520 1230
rect 968 50 1028 1230
rect 370 130 430 1150
rect 1890 130 1950 510
rect 1890 770 1950 1150
rect 770 210 830 430
rect 770 530 830 750
rect 770 850 830 1070
rect 1490 210 1550 430
rect 1490 530 1550 750
rect 1490 850 1550 1070
<< m3 >>
rect 1400 0 1600 1280
rect 680 0 880 1280
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1160 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1160 1280
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL MP2
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use PCHDL MP3
transform 1 0 1160 0 1 960
box 1160 960 2320 1280
use cut_M1M4_2x1 
transform 1 0 1400 0 1 530
box 1400 530 1600 598
use cut_M1M4_2x1 
transform 1 0 1400 0 1 690
box 1400 690 1600 758
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
use cut_M1M4_2x1 
transform 1 0 680 0 1 530
box 680 530 880 598
use cut_M1M4_2x1 
transform 1 0 680 0 1 690
box 680 690 880 758
<< labels >>
flabel locali s 1800 130 2040 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 1800 770 2040 830 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 280 450 520 510 0 FreeSans 400 0 0 0 RST
port 3 nsew
flabel locali s 680 1170 920 1230 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel m3 s 1400 0 1600 1280 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 680 0 880 1280 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
