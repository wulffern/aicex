magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1260 960
<< m1 >>
rect 90 -40 1230 40
rect 1170 40 1230 120
rect 90 120 1110 200
rect 1170 120 1230 200
rect 90 200 150 280
rect 1170 200 1230 280
rect 90 280 150 360
rect 210 280 1230 360
rect 90 360 150 440
rect 1170 360 1230 440
rect 90 440 1110 520
rect 1170 440 1230 520
rect 90 520 150 600
rect 1170 520 1230 600
rect 90 600 150 680
rect 210 600 1230 680
rect 90 680 150 760
rect 90 760 1230 840
<< m2 >>
rect 90 -40 1230 40
rect 1170 40 1230 120
rect 90 120 1110 200
rect 1170 120 1230 200
rect 90 200 150 280
rect 1170 200 1230 280
rect 90 280 150 360
rect 210 280 1230 360
rect 90 360 150 440
rect 1170 360 1230 440
rect 90 440 1110 520
rect 1170 440 1230 520
rect 90 520 150 600
rect 1170 520 1230 600
rect 90 600 150 680
rect 210 600 1230 680
rect 90 680 150 760
rect 90 760 1230 840
<< locali >>
rect 90 -40 1230 40
rect 1170 40 1230 120
rect 90 120 1110 200
rect 1170 120 1230 200
rect 90 200 150 280
rect 1170 200 1230 280
rect 90 280 150 360
rect 210 280 1230 360
rect 90 360 150 440
rect 1170 360 1230 440
rect 90 440 1110 520
rect 1170 440 1230 520
rect 90 520 150 600
rect 1170 520 1230 600
rect 90 600 150 680
rect 210 600 1230 680
rect 90 680 150 760
rect 90 760 1230 840
<< v1 >>
rect 930 -32 990 -24
rect 930 -24 990 -16
rect 930 -16 990 -8
rect 930 -8 990 0
rect 930 0 990 8
rect 930 8 990 16
rect 930 16 990 24
rect 930 24 990 32
rect 990 -32 1050 -24
rect 990 -24 1050 -16
rect 990 -16 1050 -8
rect 990 -8 1050 0
rect 990 0 1050 8
rect 990 8 1050 16
rect 990 16 1050 24
rect 990 24 1050 32
rect 1050 -32 1110 -24
rect 1050 -24 1110 -16
rect 1050 -16 1110 -8
rect 1050 -8 1110 0
rect 1050 0 1110 8
rect 1050 8 1110 16
rect 1050 16 1110 24
rect 1050 24 1110 32
rect 270 128 330 136
rect 270 136 330 144
rect 270 144 330 152
rect 270 152 330 160
rect 270 160 330 168
rect 270 168 330 176
rect 270 176 330 184
rect 270 184 330 192
rect 330 128 390 136
rect 330 136 390 144
rect 330 144 390 152
rect 330 152 390 160
rect 330 160 390 168
rect 330 168 390 176
rect 330 176 390 184
rect 330 184 390 192
rect 390 128 450 136
rect 390 136 450 144
rect 390 144 450 152
rect 390 152 450 160
rect 390 160 450 168
rect 390 168 450 176
rect 390 176 450 184
rect 390 184 450 192
rect 930 288 990 296
rect 930 296 990 304
rect 930 304 990 312
rect 930 312 990 320
rect 930 320 990 328
rect 930 328 990 336
rect 930 336 990 344
rect 930 344 990 352
rect 990 288 1050 296
rect 990 296 1050 304
rect 990 304 1050 312
rect 990 312 1050 320
rect 990 320 1050 328
rect 990 328 1050 336
rect 990 336 1050 344
rect 990 344 1050 352
rect 1050 288 1110 296
rect 1050 296 1110 304
rect 1050 304 1110 312
rect 1050 312 1110 320
rect 1050 320 1110 328
rect 1050 328 1110 336
rect 1050 336 1110 344
rect 1050 344 1110 352
rect 270 448 330 456
rect 270 456 330 464
rect 270 464 330 472
rect 270 472 330 480
rect 270 480 330 488
rect 270 488 330 496
rect 270 496 330 504
rect 270 504 330 512
rect 330 448 390 456
rect 330 456 390 464
rect 330 464 390 472
rect 330 472 390 480
rect 330 480 390 488
rect 330 488 390 496
rect 330 496 390 504
rect 330 504 390 512
rect 390 448 450 456
rect 390 456 450 464
rect 390 464 450 472
rect 390 472 450 480
rect 390 480 450 488
rect 390 488 450 496
rect 390 496 450 504
rect 390 504 450 512
rect 930 608 990 616
rect 930 616 990 624
rect 930 624 990 632
rect 930 632 990 640
rect 930 640 990 648
rect 930 648 990 656
rect 930 656 990 664
rect 930 664 990 672
rect 990 608 1050 616
rect 990 616 1050 624
rect 990 624 1050 632
rect 990 632 1050 640
rect 990 640 1050 648
rect 990 648 1050 656
rect 990 656 1050 664
rect 990 664 1050 672
rect 1050 608 1110 616
rect 1050 616 1110 624
rect 1050 624 1110 632
rect 1050 632 1110 640
rect 1050 640 1110 648
rect 1050 648 1110 656
rect 1050 656 1110 664
rect 1050 664 1110 672
rect 270 768 330 776
rect 270 776 330 784
rect 270 784 330 792
rect 270 792 330 800
rect 270 800 330 808
rect 270 808 330 816
rect 270 816 330 824
rect 270 824 330 832
rect 330 768 390 776
rect 330 776 390 784
rect 330 784 390 792
rect 330 792 390 800
rect 330 800 390 808
rect 330 808 390 816
rect 330 816 390 824
rect 330 824 390 832
rect 390 768 450 776
rect 390 776 450 784
rect 390 784 450 792
rect 390 792 450 800
rect 390 800 450 808
rect 390 808 450 816
rect 390 816 450 824
rect 390 824 450 832
<< v2 >>
rect 930 -32 990 -24
rect 930 -24 990 -16
rect 930 -16 990 -8
rect 930 -8 990 0
rect 930 0 990 8
rect 930 8 990 16
rect 930 16 990 24
rect 930 24 990 32
rect 990 -32 1050 -24
rect 990 -24 1050 -16
rect 990 -16 1050 -8
rect 990 -8 1050 0
rect 990 0 1050 8
rect 990 8 1050 16
rect 990 16 1050 24
rect 990 24 1050 32
rect 1050 -32 1110 -24
rect 1050 -24 1110 -16
rect 1050 -16 1110 -8
rect 1050 -8 1110 0
rect 1050 0 1110 8
rect 1050 8 1110 16
rect 1050 16 1110 24
rect 1050 24 1110 32
rect 270 128 330 136
rect 270 136 330 144
rect 270 144 330 152
rect 270 152 330 160
rect 270 160 330 168
rect 270 168 330 176
rect 270 176 330 184
rect 270 184 330 192
rect 330 128 390 136
rect 330 136 390 144
rect 330 144 390 152
rect 330 152 390 160
rect 330 160 390 168
rect 330 168 390 176
rect 330 176 390 184
rect 330 184 390 192
rect 390 128 450 136
rect 390 136 450 144
rect 390 144 450 152
rect 390 152 450 160
rect 390 160 450 168
rect 390 168 450 176
rect 390 176 450 184
rect 390 184 450 192
rect 930 288 990 296
rect 930 296 990 304
rect 930 304 990 312
rect 930 312 990 320
rect 930 320 990 328
rect 930 328 990 336
rect 930 336 990 344
rect 930 344 990 352
rect 990 288 1050 296
rect 990 296 1050 304
rect 990 304 1050 312
rect 990 312 1050 320
rect 990 320 1050 328
rect 990 328 1050 336
rect 990 336 1050 344
rect 990 344 1050 352
rect 1050 288 1110 296
rect 1050 296 1110 304
rect 1050 304 1110 312
rect 1050 312 1110 320
rect 1050 320 1110 328
rect 1050 328 1110 336
rect 1050 336 1110 344
rect 1050 344 1110 352
rect 270 448 330 456
rect 270 456 330 464
rect 270 464 330 472
rect 270 472 330 480
rect 270 480 330 488
rect 270 488 330 496
rect 270 496 330 504
rect 270 504 330 512
rect 330 448 390 456
rect 330 456 390 464
rect 330 464 390 472
rect 330 472 390 480
rect 330 480 390 488
rect 330 488 390 496
rect 330 496 390 504
rect 330 504 390 512
rect 390 448 450 456
rect 390 456 450 464
rect 390 464 450 472
rect 390 472 450 480
rect 390 480 450 488
rect 390 488 450 496
rect 390 496 450 504
rect 390 504 450 512
rect 930 608 990 616
rect 930 616 990 624
rect 930 624 990 632
rect 930 632 990 640
rect 930 640 990 648
rect 930 648 990 656
rect 930 656 990 664
rect 930 664 990 672
rect 990 608 1050 616
rect 990 616 1050 624
rect 990 624 1050 632
rect 990 632 1050 640
rect 990 640 1050 648
rect 990 648 1050 656
rect 990 656 1050 664
rect 990 664 1050 672
rect 1050 608 1110 616
rect 1050 616 1110 624
rect 1050 624 1110 632
rect 1050 632 1110 640
rect 1050 640 1110 648
rect 1050 648 1110 656
rect 1050 656 1110 664
rect 1050 664 1110 672
rect 270 768 330 776
rect 270 776 330 784
rect 270 784 330 792
rect 270 792 330 800
rect 270 800 330 808
rect 270 808 330 816
rect 270 816 330 824
rect 270 824 330 832
rect 330 768 390 776
rect 330 776 390 784
rect 330 784 390 792
rect 330 792 390 800
rect 330 800 390 808
rect 330 808 390 816
rect 330 816 390 824
rect 330 824 390 832
rect 390 768 450 776
rect 390 776 450 784
rect 390 784 450 792
rect 390 792 450 800
rect 390 800 450 808
rect 390 808 450 816
rect 390 816 450 824
rect 390 824 450 832
<< viali >>
rect 930 -32 990 -24
rect 930 -24 990 -16
rect 930 -16 990 -8
rect 930 -8 990 0
rect 930 0 990 8
rect 930 8 990 16
rect 930 16 990 24
rect 930 24 990 32
rect 990 -32 1050 -24
rect 990 -24 1050 -16
rect 990 -16 1050 -8
rect 990 -8 1050 0
rect 990 0 1050 8
rect 990 8 1050 16
rect 990 16 1050 24
rect 990 24 1050 32
rect 1050 -32 1110 -24
rect 1050 -24 1110 -16
rect 1050 -16 1110 -8
rect 1050 -8 1110 0
rect 1050 0 1110 8
rect 1050 8 1110 16
rect 1050 16 1110 24
rect 1050 24 1110 32
rect 270 128 330 136
rect 270 136 330 144
rect 270 144 330 152
rect 270 152 330 160
rect 270 160 330 168
rect 270 168 330 176
rect 270 176 330 184
rect 270 184 330 192
rect 330 128 390 136
rect 330 136 390 144
rect 330 144 390 152
rect 330 152 390 160
rect 330 160 390 168
rect 330 168 390 176
rect 330 176 390 184
rect 330 184 390 192
rect 390 128 450 136
rect 390 136 450 144
rect 390 144 450 152
rect 390 152 450 160
rect 390 160 450 168
rect 390 168 450 176
rect 390 176 450 184
rect 390 184 450 192
rect 930 288 990 296
rect 930 296 990 304
rect 930 304 990 312
rect 930 312 990 320
rect 930 320 990 328
rect 930 328 990 336
rect 930 336 990 344
rect 930 344 990 352
rect 990 288 1050 296
rect 990 296 1050 304
rect 990 304 1050 312
rect 990 312 1050 320
rect 990 320 1050 328
rect 990 328 1050 336
rect 990 336 1050 344
rect 990 344 1050 352
rect 1050 288 1110 296
rect 1050 296 1110 304
rect 1050 304 1110 312
rect 1050 312 1110 320
rect 1050 320 1110 328
rect 1050 328 1110 336
rect 1050 336 1110 344
rect 1050 344 1110 352
rect 270 448 330 456
rect 270 456 330 464
rect 270 464 330 472
rect 270 472 330 480
rect 270 480 330 488
rect 270 488 330 496
rect 270 496 330 504
rect 270 504 330 512
rect 330 448 390 456
rect 330 456 390 464
rect 330 464 390 472
rect 330 472 390 480
rect 330 480 390 488
rect 330 488 390 496
rect 330 496 390 504
rect 330 504 390 512
rect 390 448 450 456
rect 390 456 450 464
rect 390 464 450 472
rect 390 472 450 480
rect 390 480 450 488
rect 390 488 450 496
rect 390 496 450 504
rect 390 504 450 512
rect 930 608 990 616
rect 930 616 990 624
rect 930 624 990 632
rect 930 632 990 640
rect 930 640 990 648
rect 930 648 990 656
rect 930 656 990 664
rect 930 664 990 672
rect 990 608 1050 616
rect 990 616 1050 624
rect 990 624 1050 632
rect 990 632 1050 640
rect 990 640 1050 648
rect 990 648 1050 656
rect 990 656 1050 664
rect 990 664 1050 672
rect 1050 608 1110 616
rect 1050 616 1110 624
rect 1050 624 1110 632
rect 1050 632 1110 640
rect 1050 640 1110 648
rect 1050 648 1110 656
rect 1050 656 1110 664
rect 1050 664 1110 672
rect 270 768 330 776
rect 270 776 330 784
rect 270 784 330 792
rect 270 792 330 800
rect 270 800 330 808
rect 270 808 330 816
rect 270 816 330 824
rect 270 824 330 832
rect 330 768 390 776
rect 330 776 390 784
rect 330 784 390 792
rect 330 792 390 800
rect 330 800 390 808
rect 330 808 390 816
rect 330 816 390 824
rect 330 824 390 832
rect 390 768 450 776
rect 390 776 450 784
rect 390 784 450 792
rect 390 792 450 800
rect 390 800 450 808
rect 390 808 450 816
rect 390 816 450 824
rect 390 824 450 832
<< m3 >>
rect 90 -40 1230 40
rect 1170 40 1230 120
rect 90 120 930 200
rect 990 120 1110 200
rect 1170 120 1230 200
rect 90 200 150 280
rect 1170 200 1230 280
rect 90 280 150 360
rect 210 280 270 360
rect 330 280 1230 360
rect 90 360 150 440
rect 1170 360 1230 440
rect 90 440 1110 520
rect 1170 440 1230 520
rect 90 520 150 600
rect 1170 520 1230 600
rect 90 600 150 680
rect 210 600 1230 680
rect 90 680 150 760
rect 90 760 1230 840
<< rm3 >>
rect 930 120 990 200
rect 270 280 330 360
<< labels >>
flabel m3 s 90 -40 1230 40 0 FreeSans 400 0 0 0 B
port 1 nsew
flabel m3 s 90 760 1230 840 0 FreeSans 400 0 0 0 A
port 2 nsew
<< end >>
