magic
tech sky130A
magscale 1 2
timestamp 1660244192
<< checkpaint >>
rect 0 -768 43960 43920
<< m3 >>
rect 1548 -768 1748 13440
rect 756 -768 956 13440
<< locali >>
rect 324 498 540 558
rect 29620 10266 29836 10326
rect 756 12026 972 12086
rect 756 16026 972 16086
use SUN_PLL_KICK x1
transform 1 0 0 0 1 0
box 0 0 4056 14208
use SUN_PLL_BIAS x2
transform 1 0 0 0 1 15088
box 0 15088 4056 35280
use SUN_PLL_BUF xb1
transform 1 0 4416 0 1 176
box 4416 176 19128 12272
use SUN_PLL_LPF xb2
transform 1 0 4416 0 1 15792
box 4416 15792 43960 43920
use SUN_PLL_DIVN xh1
transform 1 0 22360 0 1 1056
box 22360 1056 37840 9420
use SUN_PLL_ROSC xh2
transform 1 0 22360 0 1 9420
box 22360 9420 28936 14828
use SUN_PLL_PFD xj1
transform 1 0 29296 0 1 9416
box 29296 9416 33352 15176
use SUN_PLL_CP xk1
transform 1 0 37672 0 1 352
box 37672 352 41728 11040
<< labels >>
flabel m3 s 1548 -768 1748 13440 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m3 s 756 -768 956 13440 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel locali s 29620 10266 29836 10326 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel locali s 756 12026 972 12086 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel locali s 756 16026 972 16086 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
