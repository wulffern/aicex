magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 50136 63000
<< locali >>
rect 49368 528 49608 62472
rect 528 528 49608 768
rect 528 62232 49608 62472
rect 528 528 768 62472
rect 49368 528 49608 62472
rect 49896 0 50136 63000
rect 0 0 50136 240
rect 0 62760 50136 63000
rect 0 0 240 63000
rect 49896 0 50136 63000
use SUN_PLL_PFD xaa0
transform 1 0 1056 0 1 1056
box 1056 1056 5112 6816
use SUN_PLL_CP xaa1
transform 1 0 5112 0 1 1056
box 5112 1056 9528 11744
use SUN_PLL_KICK xaa3
transform 1 0 9528 0 1 1056
box 9528 1056 13656 11568
use SUN_PLL_BUF xaa4
transform 1 0 13656 0 1 1056
box 13656 1056 28368 12096
use SUN_PLL_ROSC xaa5
transform 1 0 28368 0 1 1056
box 28368 1056 34944 6464
use SUN_PLL_DIVN xaa6
transform 1 0 34944 0 1 1056
box 34944 1056 49080 8092
use SUN_PLL_LPF xbb0
transform 1 0 1056 0 1 12096
box 1056 12096 40888 61944
use SUN_PLL_BIAS xbb1
transform 1 0 40888 0 1 12096
box 40888 12096 42916 30816
<< labels >>
flabel locali s 49368 528 49608 62472 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 49896 0 50136 63000 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
<< end >>
