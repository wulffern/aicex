** sch_path:
*+ /Users/wulff/pro/aicex/ip/sun_pll_sky130nm/work/../design/SUN_PLL_SKY130NM/SUN_PLL_PFD.sch
.subckt SUN_PLL_PFD CK_FB CK_REF CP_UP CP_DOWN AVDD AVSS
*.ipin CK_FB
*.ipin CK_REF
*.opin CP_UP
*.opin CP_DOWN
*.ipin AVDD
*.ipin AVSS
xa0 AVDD AVSS SUNTR_TAPCELLB_CV
xa1 CFB CK_REF CP_UP_N AVDD AVSS SUNTR_DFTSPCX1_CV
xa2 CP_UP_N CP_UP AVDD AVSS SUNTR_IVX1_CV
xa3 CP_UP_N CP_DOWN_N CFB AVDD AVSS SUNTR_NRX1_CV
xa5 CFB CK_FB CP_DOWN_N AVDD AVSS SUNTR_DFTSPCX1_CV
xa6 CP_DOWN_N CP_DOWN AVDD AVSS SUNTR_IVX1_CV
.ends
.end
