magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 1600
<< locali >>
rect 800 210 968 270
rect 800 370 968 430
rect 800 690 968 750
rect 800 1010 968 1070
rect 968 210 1028 1070
rect 1292 210 1520 270
rect 1292 370 1520 430
rect 1292 850 1520 910
rect 1292 1170 1520 1230
rect 1292 210 1352 1230
rect 370 130 430 510
rect 1920 770 2088 830
rect 1520 530 2088 590
rect 1920 1090 2088 1150
rect 1920 1410 2088 1470
rect 2088 530 2148 1470
rect 172 770 400 830
rect 172 530 800 590
rect 172 1090 400 1150
rect 172 1410 400 1470
rect 172 530 232 1470
rect 572 850 800 910
rect 572 1170 800 1230
rect 572 850 632 1230
rect 800 1490 968 1550
rect 968 1490 1520 1550
rect 968 1490 1028 1550
rect 800 1170 968 1230
rect 968 1330 1520 1390
rect 968 1170 1028 1390
rect 1520 690 1688 750
rect 1520 1010 1688 1070
rect 1688 690 1748 1070
<< m1 >>
rect 800 1330 968 1390
rect 968 1010 1520 1070
rect 968 1010 1028 1398
rect 800 530 968 590
rect 968 530 1520 590
rect 968 530 1028 598
<< poly >>
rect 280 142 2040 178
rect 280 462 2040 498
<< m3 >>
rect 1400 0 1600 1600
rect 680 0 880 1600
use NCHDL XA2
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL XA3
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL XA4a
transform 1 0 0 0 1 640
box 0 640 1160 960
use NCHDL XA4b
transform 1 0 0 0 1 960
box 0 960 1160 1280
use NCHDL XA5
transform 1 0 0 0 1 1280
box 0 1280 1160 1600
use PCHDL XB0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL XB1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL XB3a
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use PCHDL XB3b
transform 1 0 1160 0 1 960
box 1160 960 2320 1280
use PCHDL XB4
transform 1 0 1160 0 1 1280
box 1160 1280 2320 1600
use cut_M1M2_2x1 
transform 1 0 680 0 1 1330
box 680 1330 880 1398
use cut_M1M2_2x1 
transform 1 0 1400 0 1 1010
box 1400 1010 1600 1078
use cut_M1M2_2x1 
transform 1 0 680 0 1 530
box 680 530 880 598
use cut_M1M2_2x1 
transform 1 0 1400 0 1 530
box 1400 530 1600 598
use cut_M1M4_2x1 
transform 1 0 1400 0 1 50
box 1400 50 1600 118
use cut_M1M4_2x1 
transform 1 0 1400 0 1 1330
box 1400 1330 1600 1398
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
use cut_M1M4_2x1 
transform 1 0 680 0 1 1330
box 680 1330 880 1398
<< labels >>
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 680 1490 920 1550 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel m3 s 1400 0 1600 1600 0 FreeSans 400 0 0 0 AVDD
port 3 nsew
flabel m3 s 680 0 880 1600 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
<< end >>
