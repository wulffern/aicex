magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 11280 4800
<< m3 >>
rect 12 760 5680 820
rect 12 1720 5680 1780
rect 12 2680 5680 2740
rect 12 3640 5680 3700
rect 12 4600 5680 4660
rect 12 760 72 4660
rect 5680 -40 11288 20
rect 5680 920 11288 980
rect 5680 1880 11288 1940
rect 5680 2840 11288 2900
rect 5680 3800 11288 3860
rect 11288 -40 11348 3860
use CAP_BSSW_CV XCAPB0
transform 1 0 0 0 1 0
box 0 0 11280 960
use CAP_BSSW_CV XCAPB1
transform 1 0 0 0 1 960
box 0 960 11280 1920
use CAP_BSSW_CV XCAPB2
transform 1 0 0 0 1 1920
box 0 1920 11280 2880
use CAP_BSSW_CV XCAPB3
transform 1 0 0 0 1 2880
box 0 2880 11280 3840
use CAP_BSSW_CV XCAPB4
transform 1 0 0 0 1 3840
box 0 3840 11280 4800
<< labels >>
flabel m3 s 120 2680 11240 2760 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel m3 s 120 -40 11240 40 0 FreeSans 400 0 0 0 B
port 2 nsew
<< end >>
