magic
tech sky130A
magscale 1 2
timestamp 1660083337
<< checkpaint >>
rect 0 0 648 2860
<< ppolyres >>
rect 162 -110 270 110
rect 378 -110 486 110
rect 162 110 270 330
rect 378 110 486 330
rect 162 330 270 550
rect 378 330 486 550
rect 162 550 270 770
rect 378 550 486 770
rect 162 770 270 990
rect 378 770 486 990
rect 162 990 270 1210
rect 378 990 486 1210
rect 162 1210 270 1430
rect 378 1210 486 1430
rect 162 1430 270 1650
rect 378 1430 486 1650
rect 162 1650 270 1870
rect 378 1650 486 1870
rect 162 1870 270 2090
rect 378 1870 486 2090
rect 162 2090 270 2310
rect 378 2090 486 2310
rect 162 2310 270 2530
rect 378 2310 486 2530
<< poly >>
rect -54 -110 54 110
rect 594 -110 702 110
rect -54 110 54 330
rect 594 110 702 330
rect -54 330 54 550
rect 594 330 702 550
rect -54 550 54 770
rect 594 550 702 770
rect -54 770 54 990
rect 594 770 702 990
rect -54 990 54 1210
rect 594 990 702 1210
rect -54 1210 54 1430
rect 594 1210 702 1430
rect -54 1430 54 1650
rect 594 1430 702 1650
rect -54 1650 54 1870
rect 594 1650 702 1870
rect -54 1870 54 2090
rect 594 1870 702 2090
rect -54 2090 54 2310
rect 594 2090 702 2310
rect -54 2310 54 2530
rect 594 2310 702 2530
<< xpolycontact >>
rect 162 -110 270 110
rect 378 -110 486 110
rect 162 110 270 330
rect 378 110 486 330
rect 162 2090 270 2310
rect 378 2090 486 2310
rect 162 2310 270 2530
rect 378 2310 486 2530
<< locali >>
rect 162 -110 486 110
rect 162 110 486 330
rect 162 2090 270 2310
rect 378 2090 486 2310
rect 162 2310 270 2530
rect 378 2310 486 2530
rect 162 2530 270 2750
rect 378 2530 486 2750
rect -54 2750 270 2970
rect -54 2750 270 2970
rect 378 2750 702 2970
rect 378 2750 702 2970
<< pwell >>
rect -54 -110 702 2970
<< labels >>
flabel locali s -54 2750 270 2970 0 FreeSans 400 0 0 0 N
port 1 nsew
flabel locali s 378 2750 702 2970 0 FreeSans 400 0 0 0 P
port 2 nsew
<< end >>
