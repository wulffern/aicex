magic
tech sky130A
magscale 1 2
timestamp 1660660914
<< checkpaint >>
rect -1440 -1644 14040 6720
<< locali >>
rect 0 -204 12600 -144
rect 0 -204 12600 -144
rect 13120 -924 13320 6000
rect -720 -924 13320 -724
rect -720 5800 13320 6000
rect -720 -924 -520 6000
rect 13120 -924 13320 6000
rect 13840 -1644 14040 6720
rect -1440 -1644 14040 -1444
rect -1440 6520 14040 6720
rect -1440 -1644 -1240 6720
rect 13840 -1644 14040 6720
rect 756 5162 972 5222
rect 10404 498 10620 558
<< m3 >>
rect 394 -204 470 4078
rect 4570 -204 4646 4078
rect 5434 -204 5510 4078
rect 9610 -204 9686 4078
rect 10474 -204 10550 4078
rect 756 -924 956 5280
rect 4084 -924 4284 5280
rect 5796 -924 5996 5280
rect 9124 -924 9324 5280
rect 10836 -924 11036 5280
rect 1548 -1644 1748 5280
rect 3292 -1644 3492 5280
rect 6588 -1644 6788 5280
rect 8332 -1644 8532 5280
rect 11628 -1644 11828 5280
<< m2 >>
rect 4608 498 4988 574
rect 4988 5238 5856 5314
rect 4988 498 5064 5314
rect 5796 5162 5904 5238
rect 9648 498 10028 574
rect 10028 5238 10896 5314
rect 10028 498 10104 5314
rect 10836 5162 10944 5238
rect 480 574 2468 650
rect 2468 5238 4128 5314
rect 2468 498 2544 5314
rect 432 498 540 574
rect 4068 5162 4176 5238
rect 5520 574 7508 650
rect 7508 5238 9168 5314
rect 7508 498 7584 5314
rect 5472 498 5580 574
rect 9108 5162 9216 5238
rect 184 5074 432 5150
rect 184 1554 432 1630
rect 184 1554 260 5150
rect 4608 5074 4780 5150
rect 4608 1554 4780 1630
rect 4780 1554 4856 5150
rect 5224 5074 5472 5150
rect 5224 1554 5472 1630
rect 5224 1554 5300 5150
rect 9648 5074 9820 5150
rect 9648 1554 9820 1630
rect 9820 1554 9896 5150
rect 10264 5074 10512 5150
rect 10264 1554 10512 1630
rect 10264 1554 10340 5150
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xc0
transform 1 0 0 0 1 0
box 0 0 2520 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xd0
transform -1 0 5040 0 1 0
box 5040 0 7560 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xe0
transform 1 0 5040 0 1 0
box 5040 0 7560 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xf0
transform -1 0 10080 0 1 0
box 10080 0 12600 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xg0
transform 1 0 10080 0 1 0
box 10080 0 12600 5280
use cut_M1M4_2x1 
transform 1 0 332 0 1 4018
box 332 4018 532 4094
use cut_M1M4_2x1 
transform 1 0 332 0 1 -204
box 332 -204 532 -128
use cut_M1M4_2x1 
transform 1 0 4508 0 1 4018
box 4508 4018 4708 4094
use cut_M1M4_2x1 
transform 1 0 4508 0 1 -204
box 4508 -204 4708 -128
use cut_M1M4_2x1 
transform 1 0 5372 0 1 4018
box 5372 4018 5572 4094
use cut_M1M4_2x1 
transform 1 0 5372 0 1 -204
box 5372 -204 5572 -128
use cut_M1M4_2x1 
transform 1 0 9548 0 1 4018
box 9548 4018 9748 4094
use cut_M1M4_2x1 
transform 1 0 9548 0 1 -204
box 9548 -204 9748 -128
use cut_M1M4_2x1 
transform 1 0 10412 0 1 4018
box 10412 4018 10612 4094
use cut_M1M4_2x1 
transform 1 0 10412 0 1 -204
box 10412 -204 10612 -128
use cut_M1M4_2x2 
transform 1 0 756 0 1 -924
box 756 -924 956 -724
use cut_M1M4_2x2 
transform 1 0 4084 0 1 -924
box 4084 -924 4284 -724
use cut_M1M4_2x2 
transform 1 0 5796 0 1 -924
box 5796 -924 5996 -724
use cut_M1M4_2x2 
transform 1 0 9124 0 1 -924
box 9124 -924 9324 -724
use cut_M1M4_2x2 
transform 1 0 10836 0 1 -924
box 10836 -924 11036 -724
use cut_M1M4_2x2 
transform 1 0 1548 0 1 -1644
box 1548 -1644 1748 -1444
use cut_M1M4_2x2 
transform 1 0 3292 0 1 -1644
box 3292 -1644 3492 -1444
use cut_M1M4_2x2 
transform 1 0 6588 0 1 -1644
box 6588 -1644 6788 -1444
use cut_M1M4_2x2 
transform 1 0 8332 0 1 -1644
box 8332 -1644 8532 -1444
use cut_M1M4_2x2 
transform 1 0 11628 0 1 -1644
box 11628 -1644 11828 -1444
use cut_M1M3_2x1 
transform 1 0 4500 0 1 498
box 4500 498 4700 574
use cut_M1M3_2x1 
transform 1 0 5796 0 1 5162
box 5796 5162 5996 5238
use cut_M1M3_2x1 
transform 1 0 9540 0 1 498
box 9540 498 9740 574
use cut_M1M3_2x1 
transform 1 0 10836 0 1 5162
box 10836 5162 11036 5238
use cut_M1M3_2x1 
transform 1 0 324 0 1 498
box 324 498 524 574
use cut_M1M3_2x1 
transform 1 0 4068 0 1 5162
box 4068 5162 4268 5238
use cut_M1M3_2x1 
transform 1 0 5364 0 1 498
box 5364 498 5564 574
use cut_M1M3_2x1 
transform 1 0 9108 0 1 5162
box 9108 5162 9308 5238
use cut_M1M3_2x1 
transform 1 0 340 0 1 5074
box 340 5074 540 5150
use cut_M1M3_2x1 
transform 1 0 340 0 1 1554
box 340 1554 540 1630
use cut_M1M3_2x1 
transform 1 0 4500 0 1 5074
box 4500 5074 4700 5150
use cut_M1M3_2x1 
transform 1 0 4500 0 1 1554
box 4500 1554 4700 1630
use cut_M1M3_2x1 
transform 1 0 5380 0 1 5074
box 5380 5074 5580 5150
use cut_M1M3_2x1 
transform 1 0 5380 0 1 1554
box 5380 1554 5580 1630
use cut_M1M3_2x1 
transform 1 0 9540 0 1 5074
box 9540 5074 9740 5150
use cut_M1M3_2x1 
transform 1 0 9540 0 1 1554
box 9540 1554 9740 1630
use cut_M1M3_2x1 
transform 1 0 10420 0 1 5074
box 10420 5074 10620 5150
use cut_M1M3_2x1 
transform 1 0 10420 0 1 1554
box 10420 1554 10620 1630
<< labels >>
flabel locali s 0 -204 12600 -144 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew
flabel locali s 13120 -924 13320 6000 0 FreeSans 400 0 0 0 AVSS
port 5 nsew
flabel locali s 13840 -1644 14040 6720 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 756 5162 972 5222 0 FreeSans 400 0 0 0 CK_FB
port 2 nsew
flabel locali s 10404 498 10620 558 0 FreeSans 400 0 0 0 CK
port 3 nsew
<< end >>
