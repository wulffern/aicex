magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 14080
<< locali >>
rect 1380 4530 1534 4590
rect 1534 8770 1740 8830
rect 1534 6210 1740 6270
rect 1534 4530 1594 8830
rect 146 2370 360 2430
rect 146 2690 360 2750
rect 146 7490 360 7550
rect 146 11650 360 11710
rect 146 2370 206 11710
rect 360 11650 514 11710
rect 514 12050 720 12110
rect 514 11650 574 12110
rect 506 13170 720 13230
rect 360 12290 506 12350
rect 506 12290 566 13230
rect 1380 13650 1534 13710
rect 1534 12610 1740 12670
rect 1534 12610 1594 13710
rect 506 4050 720 4110
rect 506 8850 720 8910
rect 506 4050 566 8910
rect 270 12930 450 12990
rect 270 13570 450 13630
rect 270 13250 450 13310
rect 630 6290 810 6350
rect 630 5010 810 5070
rect 270 2050 450 2110
rect 270 9090 450 9150
<< m1 >>
rect 1380 8690 1534 8750
rect 1534 4290 1740 4350
rect 1534 4930 1740 4990
rect 1534 4290 1594 8758
rect 360 2050 514 2110
rect 360 3010 514 3070
rect 514 2050 574 3078
rect 360 9090 514 9150
rect 360 10050 514 10110
rect 514 9090 574 10118
rect 146 450 360 510
rect 146 9730 360 9790
rect 146 11970 360 12030
rect 146 450 206 12038
rect 360 11970 514 12030
rect 514 12690 720 12750
rect 514 11970 574 12758
<< m3 >>
rect 1290 0 1474 14080
rect 630 0 814 14080
rect 1290 0 1474 14080
rect 630 0 814 14080
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use TAPCELLB_CV XA0
transform 1 0 0 0 1 0
box 0 0 2100 320
use SARKICKHX1_CV XA1
transform 1 0 0 0 1 320
box 0 320 2100 2560
use SARCMPHX1_CV XA2
transform 1 0 0 0 1 2560
box 0 2560 2100 4800
use IVX4_CV XA2a
transform 1 0 0 0 1 4800
box 0 4800 2100 6080
use IVX4_CV XA3a
transform 1 0 0 0 1 6080
box 0 6080 2100 7360
use SARCMPHX1_CV XA3
transform 1 0 0 0 1 7360
box 0 7360 2100 9600
use SARKICKHX1_CV XA4
transform 1 0 0 0 1 9600
box 0 9600 2100 11840
use IVX1_CV XA9
transform 1 0 0 0 1 11840
box 0 11840 2100 12160
use NDX1_CV XA10
transform 1 0 0 0 1 12160
box 0 12160 2100 12800
use NRX1_CV XA11
transform 1 0 0 0 1 12800
box 0 12800 2100 13440
use IVX1_CV XA12
transform 1 0 0 0 1 13440
box 0 13440 2100 13760
use TAPCELLB_CV XA13
transform 1 0 0 0 1 13760
box 0 13760 2100 14080
use DMY_CV XA14
transform 1 0 0 0 1 14080
box 0 14080 0 14080
use cut_M1M2_2x1 
transform 1 0 1290 0 1 8690
box 1290 8690 1474 8758
use cut_M1M2_2x1 
transform 1 0 1650 0 1 4290
box 1650 4290 1834 4358
use cut_M1M2_2x1 
transform 1 0 1650 0 1 4930
box 1650 4930 1834 4998
use cut_M1M2_2x1 
transform 1 0 266 0 1 2050
box 266 2050 450 2118
use cut_M1M2_2x1 
transform 1 0 266 0 1 3010
box 266 3010 450 3078
use cut_M1M2_2x1 
transform 1 0 266 0 1 9090
box 266 9090 450 9158
use cut_M1M2_2x1 
transform 1 0 266 0 1 10050
box 266 10050 450 10118
use cut_M1M2_2x1 
transform 1 0 270 0 1 450
box 270 450 454 518
use cut_M1M2_2x1 
transform 1 0 270 0 1 9730
box 270 9730 454 9798
use cut_M1M2_2x1 
transform 1 0 270 0 1 11970
box 270 11970 454 12038
use cut_M1M2_2x1 
transform 1 0 270 0 1 11970
box 270 11970 454 12038
use cut_M1M2_2x1 
transform 1 0 630 0 1 12690
box 630 12690 814 12758
<< labels >>
flabel locali s 270 12930 450 12990 0 FreeSans 400 0 0 0 CK_SAMPLE
port 1 nsew
flabel locali s 270 13570 450 13630 0 FreeSans 400 0 0 0 CK_CMP
port 2 nsew
flabel locali s 270 13250 450 13310 0 FreeSans 400 0 0 0 DONE
port 3 nsew
flabel locali s 630 6290 810 6350 0 FreeSans 400 0 0 0 CNO
port 4 nsew
flabel locali s 630 5010 810 5070 0 FreeSans 400 0 0 0 CPO
port 5 nsew
flabel locali s 270 2050 450 2110 0 FreeSans 400 0 0 0 CPI
port 6 nsew
flabel locali s 270 9090 450 9150 0 FreeSans 400 0 0 0 CNI
port 7 nsew
flabel m3 s 1290 0 1474 14080 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 14080 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
