magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 13120
<< locali >>
rect 360 5250 498 5310
rect 498 4050 720 4110
rect 498 4050 558 5310
rect 360 7810 498 7870
rect 498 6610 720 6670
rect 498 6610 558 7870
rect 1422 3970 1620 4030
rect 1260 3730 1422 3790
rect 1422 3730 1482 4030
rect 360 10690 498 10750
rect 498 10450 720 10510
rect 498 10450 558 10750
rect 330 10690 390 11070
rect 390 11590 498 11650
rect 498 11410 720 11470
rect 498 11410 558 11650
rect 390 11650 450 11710
rect 390 11910 498 11970
rect 498 11730 720 11790
rect 498 11730 558 11970
rect 390 11970 450 12030
rect 360 12610 498 12670
rect 498 12210 720 12270
rect 498 12210 558 12670
rect 1260 7890 1398 7950
rect 1398 9090 1620 9150
rect 1398 7890 1458 9150
<< m1 >>
rect 360 6530 498 6590
rect 498 2770 720 2830
rect 498 2770 558 6598
rect 1620 10370 1758 10430
rect 1260 690 1758 750
rect 1758 690 1818 10438
rect 360 11330 498 11390
rect 498 10130 720 10190
rect 498 10130 558 11398
rect 1260 5330 1398 5390
rect 1398 9730 1620 9790
rect 1398 5330 1458 9798
<< m3 >>
rect 1712 4370 1772 8394
rect 1170 0 1354 13120
rect 630 0 814 13120
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use SARMRYX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 1980 3840
use SWX4_CV XA2
transform 1 0 0 0 1 3840
box 0 3840 1980 5120
use SWX4_CV XA3
transform 1 0 0 0 1 5120
box 0 5120 1980 6400
use SWX4_CV XA4
transform 1 0 0 0 1 6400
box 0 6400 1980 7680
use SWX4_CV XA5
transform 1 0 0 0 1 7680
box 0 7680 1980 8960
use SARCEX1_CV XA6
transform 1 0 0 0 1 8960
box 0 8960 1980 10240
use IVX1_CV XA7
transform 1 0 0 0 1 10240
box 0 10240 1980 10560
use IVX1_CV XA8
transform 1 0 0 0 1 10560
box 0 10560 1980 10880
use NDX1_CV XA9
transform 1 0 0 0 1 10880
box 0 10880 1980 11520
use IVX1_CV XA10
transform 1 0 0 0 1 11520
box 0 11520 1980 11840
use NRX1_CV XA11
transform 1 0 0 0 1 11840
box 0 11840 1980 12480
use IVX1_CV XA12
transform 1 0 0 0 1 12480
box 0 12480 1980 12800
use TAPCELLB_CV XA13
transform 1 0 0 0 1 12800
box 0 12800 1980 13120
use DMY_CV XA14
transform 1 0 0 0 1 13120
box 0 13120 0 13120
use cut_M1M2_2x1 
transform 1 0 270 0 1 6530
box 270 6530 454 6598
use cut_M1M2_2x1 
transform 1 0 630 0 1 2770
box 630 2770 814 2838
use cut_M1M2_2x1 
transform 1 0 1530 0 1 10370
box 1530 10370 1714 10438
use cut_M1M2_2x1 
transform 1 0 1170 0 1 690
box 1170 690 1354 758
use cut_M1M2_2x1 
transform 1 0 270 0 1 11330
box 270 11330 454 11398
use cut_M1M2_2x1 
transform 1 0 630 0 1 10130
box 630 10130 814 10198
use cut_M1M2_2x1 
transform 1 0 1170 0 1 5330
box 1170 5330 1354 5398
use cut_M1M2_2x1 
transform 1 0 1530 0 1 9730
box 1530 9730 1714 9798
use cut_M1M4_2x1 
transform 1 0 266 0 1 5246
box 266 5246 450 5314
use cut_M1M4_1x2 
transform 1 0 946 0 1 5268
box 946 5268 1014 5452
use cut_M1M4_1x2 
transform 1 0 1082 0 1 6548
box 1082 6548 1150 6732
use cut_M1M4_1x2 
transform 1 0 1218 0 1 7828
box 1218 7828 1286 8012
use cut_M2M3_2x1 
transform 1 0 1166 0 1 686
box 1166 686 1350 754
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
<< labels >>
flabel m2 s 266 2046 450 2114 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1530 3650 1710 3710 0 FreeSans 400 0 0 0 RST_N
port 2 nsew
flabel m2 s 266 446 450 514 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 270 3010 450 3070 0 FreeSans 400 0 0 0 CMP_ON
port 4 nsew
flabel m2 s 1166 686 1350 754 0 FreeSans 400 0 0 0 ENO
port 5 nsew
flabel m3 s 266 5246 450 5314 0 FreeSans 400 0 0 0 CN1
port 6 nsew
flabel m3 s 946 5268 1014 5452 0 FreeSans 400 0 0 0 CP1
port 7 nsew
flabel m3 s 1082 6548 1150 6732 0 FreeSans 400 0 0 0 CP0
port 8 nsew
flabel m3 s 1218 7828 1286 8012 0 FreeSans 400 0 0 0 CN0
port 9 nsew
flabel locali s 270 12290 450 12350 0 FreeSans 400 0 0 0 CEIN
port 10 nsew
flabel locali s 1170 12690 1350 12750 0 FreeSans 400 0 0 0 CEO
port 11 nsew
flabel locali s 270 9410 450 9470 0 FreeSans 400 0 0 0 CKS
port 12 nsew
flabel locali s 630 10770 810 10830 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 1650 4370 1834 4554 0 FreeSans 400 0 0 0 VREF
port 14 nsew
flabel m3 s 1170 0 1354 13120 0 FreeSans 400 0 0 0 AVDD
port 15 nsew
flabel m3 s 630 0 814 13120 0 FreeSans 400 0 0 0 AVSS
port 16 nsew
<< end >>
