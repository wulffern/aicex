magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 1280
<< locali >>
rect 1490 530 1550 750
rect 1490 850 1550 1070
rect 800 210 968 270
rect 800 530 968 590
rect 800 690 968 750
rect 968 210 1028 750
rect 1292 370 1520 430
rect 800 1170 1292 1230
rect 1292 370 1352 1230
rect 1520 50 1688 110
rect 1688 1090 1920 1150
rect 1688 50 1748 1150
rect 680 50 1640 110
<< poly >>
rect 280 462 2040 498
rect 280 782 2040 818
rect 280 1102 2040 1138
<< m3 >>
rect 1400 0 1600 1280
rect 680 0 880 1280
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1160 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1160 1280
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL MP2
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use PCHDL MP3
transform 1 0 1160 0 1 960
box 1160 960 2320 1280
use cut_M1M4_2x1 
transform 1 0 1400 0 1 210
box 1400 210 1600 278
use cut_M1M4_2x1 
transform 1 0 1400 0 1 1170
box 1400 1170 1600 1238
use cut_M1M4_2x1 
transform 1 0 680 0 1 370
box 680 370 880 438
use cut_M1M4_2x1 
transform 1 0 680 0 1 850
box 680 850 880 918
use cut_M1M4_2x1 
transform 1 0 680 0 1 1010
box 680 1010 880 1078
<< labels >>
flabel locali s 2200 120 2440 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -120 120 120 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 280 770 520 830 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel locali s 280 450 520 510 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 1800 130 2040 190 0 FreeSans 400 0 0 0 RST_N
port 5 nsew
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 EN
port 6 nsew
flabel locali s 1400 370 1640 430 0 FreeSans 400 0 0 0 ENO
port 7 nsew
flabel m3 s 1400 0 1600 1280 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 680 0 880 1280 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
