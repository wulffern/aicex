magic
tech sky130A
magscale 1 2
timestamp 1659304800
<< checkpaint >>
rect 0 0 1928 4140
<< locali >>
rect 0 0 1928 112
rect 0 0 1928 112
rect 0 0 112 4140
rect 0 4028 1928 4140
rect 1816 0 1928 4140
rect 0 0 1928 112
rect 1018 3390 1342 3610
rect 586 3390 910 3610
<< ptapc >>
rect 4 0 84 80
rect 84 0 164 80
rect 164 0 244 80
rect 244 0 324 80
rect 324 0 404 80
rect 404 0 484 80
rect 484 0 564 80
rect 564 0 644 80
rect 644 0 724 80
rect 724 0 804 80
rect 804 0 884 80
rect 884 0 964 80
rect 964 0 1044 80
rect 1044 0 1124 80
rect 1124 0 1204 80
rect 1204 0 1284 80
rect 1284 0 1364 80
rect 1364 0 1444 80
rect 1444 0 1524 80
rect 1524 0 1604 80
rect 1604 0 1684 80
rect 1684 0 1764 80
rect 1764 0 1844 80
rect 1844 0 1924 80
rect 0 30 80 110
rect 0 110 80 190
rect 0 190 80 270
rect 0 270 80 350
rect 0 350 80 430
rect 0 430 80 510
rect 0 510 80 590
rect 0 590 80 670
rect 0 670 80 750
rect 0 750 80 830
rect 0 830 80 910
rect 0 910 80 990
rect 0 990 80 1070
rect 0 1070 80 1150
rect 0 1150 80 1230
rect 0 1230 80 1310
rect 0 1310 80 1390
rect 0 1390 80 1470
rect 0 1470 80 1550
rect 0 1550 80 1630
rect 0 1630 80 1710
rect 0 1710 80 1790
rect 0 1790 80 1870
rect 0 1870 80 1950
rect 0 1950 80 2030
rect 0 2030 80 2110
rect 0 2110 80 2190
rect 0 2190 80 2270
rect 0 2270 80 2350
rect 0 2350 80 2430
rect 0 2430 80 2510
rect 0 2510 80 2590
rect 0 2590 80 2670
rect 0 2670 80 2750
rect 0 2750 80 2830
rect 0 2830 80 2910
rect 0 2910 80 2990
rect 0 2990 80 3070
rect 0 3070 80 3150
rect 0 3150 80 3230
rect 0 3230 80 3310
rect 0 3310 80 3390
rect 0 3390 80 3470
rect 0 3470 80 3550
rect 0 3550 80 3630
rect 0 3630 80 3710
rect 0 3710 80 3790
rect 0 3790 80 3870
rect 0 3870 80 3950
rect 0 3950 80 4030
rect 0 4030 80 4110
rect 4 4028 84 4108
rect 84 4028 164 4108
rect 164 4028 244 4108
rect 244 4028 324 4108
rect 324 4028 404 4108
rect 404 4028 484 4108
rect 484 4028 564 4108
rect 564 4028 644 4108
rect 644 4028 724 4108
rect 724 4028 804 4108
rect 804 4028 884 4108
rect 884 4028 964 4108
rect 964 4028 1044 4108
rect 1044 4028 1124 4108
rect 1124 4028 1204 4108
rect 1204 4028 1284 4108
rect 1284 4028 1364 4108
rect 1364 4028 1444 4108
rect 1444 4028 1524 4108
rect 1524 4028 1604 4108
rect 1604 4028 1684 4108
rect 1684 4028 1764 4108
rect 1764 4028 1844 4108
rect 1844 4028 1924 4108
rect 1816 30 1896 110
rect 1816 110 1896 190
rect 1816 190 1896 270
rect 1816 270 1896 350
rect 1816 350 1896 430
rect 1816 430 1896 510
rect 1816 510 1896 590
rect 1816 590 1896 670
rect 1816 670 1896 750
rect 1816 750 1896 830
rect 1816 830 1896 910
rect 1816 910 1896 990
rect 1816 990 1896 1070
rect 1816 1070 1896 1150
rect 1816 1150 1896 1230
rect 1816 1230 1896 1310
rect 1816 1310 1896 1390
rect 1816 1390 1896 1470
rect 1816 1470 1896 1550
rect 1816 1550 1896 1630
rect 1816 1630 1896 1710
rect 1816 1710 1896 1790
rect 1816 1790 1896 1870
rect 1816 1870 1896 1950
rect 1816 1950 1896 2030
rect 1816 2030 1896 2110
rect 1816 2110 1896 2190
rect 1816 2190 1896 2270
rect 1816 2270 1896 2350
rect 1816 2350 1896 2430
rect 1816 2430 1896 2510
rect 1816 2510 1896 2590
rect 1816 2590 1896 2670
rect 1816 2670 1896 2750
rect 1816 2750 1896 2830
rect 1816 2830 1896 2910
rect 1816 2910 1896 2990
rect 1816 2990 1896 3070
rect 1816 3070 1896 3150
rect 1816 3150 1896 3230
rect 1816 3230 1896 3310
rect 1816 3310 1896 3390
rect 1816 3390 1896 3470
rect 1816 3470 1896 3550
rect 1816 3550 1896 3630
rect 1816 3630 1896 3710
rect 1816 3710 1896 3790
rect 1816 3790 1896 3870
rect 1816 3870 1896 3950
rect 1816 3950 1896 4030
rect 1816 4030 1896 4110
<< ptap >>
rect 0 0 1928 112
rect 0 0 112 4140
rect 0 4028 1928 4140
rect 1816 0 1928 4140
use SUNTR_RES12 XA1
transform 1 0 640 0 1 640
box 640 640 1288 3500
<< labels >>
flabel locali s 0 0 1928 112 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 1018 3390 1342 3610 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 586 3390 910 3610 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
