magic
tech sky130A
magscale 1 2
timestamp 1661026409
<< checkpaint >>
rect 0 0 4056 14208
<< m3 >>
rect 1524 0 1724 14208
rect 1516 384 1732 1120
rect 1516 384 1732 1472
rect 1516 384 1732 1824
rect 1516 384 1732 4640
rect 2316 0 2516 14208
rect 2308 0 2524 1120
rect 2308 0 2524 1472
rect 2308 0 2524 1824
rect 2308 0 2524 4640
rect 2316 0 2516 14208
rect 1524 0 1724 14208
<< locali >>
rect 384 384 3672 624
rect 384 13584 3672 13824
rect 384 384 624 13824
rect 3432 384 3672 13824
rect 0 0 4056 240
rect 0 13968 4056 14208
rect 0 0 240 14208
rect 3816 0 4056 14208
rect 1404 1766 1584 1826
rect 1200 1970 1404 2030
rect 1200 4786 1404 4846
rect 1404 1766 1464 4846
rect 1524 1706 1632 1766
rect 1404 4934 1584 4994
rect 1200 5138 1404 5198
rect 1404 4934 1464 5198
rect 1524 4874 1632 4934
rect 1404 5286 1584 5346
rect 1200 5490 1404 5550
rect 1200 8306 1404 8366
rect 1404 5286 1464 8366
rect 1524 5226 1632 5286
rect 1404 8454 1584 8514
rect 1200 8658 1404 8718
rect 1404 8454 1464 8718
rect 1524 8394 1632 8454
rect 1404 8806 1584 8866
rect 1200 9010 1404 9070
rect 1200 11826 1404 11886
rect 1404 8806 1464 11886
rect 1524 8746 1632 8806
rect 1404 11974 1584 12034
rect 1200 12178 1404 12238
rect 1404 11974 1464 12238
rect 1524 11914 1632 11974
rect 1404 12326 1584 12386
rect 1200 12882 1404 12942
rect 1404 12326 1464 12942
rect 1524 12266 1632 12326
rect 1524 12794 1740 12854
rect 1524 13322 1740 13382
rect 1092 1266 1308 1326
rect 1524 1354 1740 1414
<< m1 >>
rect 1200 13234 1368 13294
rect 1368 12794 1632 12854
rect 1368 12794 1428 13302
rect 972 1618 1200 1678
rect 972 1354 1632 1414
rect 972 12530 1200 12590
rect 972 1354 1032 12598
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV xa1a0
transform 1 0 768 0 1 768
box 768 768 3288 1120
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa1b0
transform 1 0 768 0 1 1120
box 768 1120 3288 1472
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa1c0
transform 1 0 768 0 1 1472
box 768 1472 3288 1824
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX8_CV xa1d0
transform 1 0 768 0 1 1824
box 768 1824 3288 4640
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa20
transform 1 0 768 0 1 4640
box 768 4640 3288 4992
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa3a0
transform 1 0 768 0 1 4992
box 768 4992 3288 5344
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX8_CV xa3b0
transform 1 0 768 0 1 5344
box 768 5344 3288 8160
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa40
transform 1 0 768 0 1 8160
box 768 8160 3288 8512
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa5a0
transform 1 0 768 0 1 8512
box 768 8512 3288 8864
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX8_CV xa5b0
transform 1 0 768 0 1 8864
box 768 8864 3288 11680
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa60
transform 1 0 768 0 1 11680
box 768 11680 3288 12032
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa70
transform 1 0 768 0 1 12032
box 768 12032 3288 12384
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NRX1_CV xa80
transform 1 0 768 0 1 12384
box 768 12384 3288 13088
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa90
transform 1 0 768 0 1 13088
box 768 13088 3288 13440
use cut_M1M4_2x1 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 
transform 1 0 2316 0 1 0
box 2316 0 2516 76
use cut_M1M4_2x1 
transform 1 0 2316 0 1 0
box 2316 0 2516 76
use cut_M1M4_2x1 
transform 1 0 2316 0 1 0
box 2316 0 2516 76
use cut_M1M4_2x1 
transform 1 0 2316 0 1 0
box 2316 0 2516 76
use cut_M1M2_2x1 
transform 1 0 1092 0 1 13234
box 1092 13234 1276 13302
use cut_M1M2_2x1 
transform 1 0 1524 0 1 12794
box 1524 12794 1708 12862
use cut_M1M2_2x1 
transform 1 0 1092 0 1 1618
box 1092 1618 1276 1686
use cut_M1M2_2x1 
transform 1 0 1524 0 1 1354
box 1524 1354 1708 1422
use cut_M1M2_2x1 
transform 1 0 1092 0 1 12530
box 1092 12530 1276 12598
<< labels >>
flabel m3 s 1524 0 1724 14208 0 FreeSans 400 0 0 0 AVSS
port 5 nsew
flabel m3 s 2316 0 2516 14208 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 1524 12794 1740 12854 0 FreeSans 400 0 0 0 KICK
port 2 nsew
flabel locali s 1524 13322 1740 13382 0 FreeSans 400 0 0 0 KICK_N
port 3 nsew
flabel locali s 1092 1266 1308 1326 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew
flabel locali s 1524 1354 1740 1414 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 6 nsew
<< end >>
