magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 30 8976 1574
<< m1 >>
rect 2308 380 2376 1604
rect 6796 0 6864 1224
rect 2572 0 2640 540
rect 2572 836 2640 1604
rect 6532 0 6600 540
rect 6532 836 6600 1604
rect 2044 0 2112 996
rect 2044 1292 2112 1604
rect 2836 0 2904 996
rect 2836 1292 2904 1604
rect 6268 0 6336 996
rect 6268 1292 6336 1604
rect 7060 0 7128 996
rect 7060 1292 7128 1604
rect 1516 0 1584 768
rect 1516 1064 1584 1604
rect 1780 0 1848 768
rect 1780 1064 1848 1604
rect 3100 0 3168 768
rect 3100 1064 3168 1604
rect 3364 0 3432 768
rect 3364 1064 3432 1604
rect 5740 0 5808 768
rect 5740 1064 5808 1604
rect 6004 0 6072 768
rect 6004 1064 6072 1604
rect 7324 0 7392 768
rect 7324 1064 7392 1604
rect 7588 0 7656 768
rect 7588 1064 7656 1604
rect 460 0 528 312
rect 460 608 528 1604
rect 724 0 792 312
rect 724 608 792 1604
rect 988 0 1056 312
rect 988 608 1056 1604
rect 1252 0 1320 312
rect 1252 608 1320 1604
rect 3628 0 3696 312
rect 3628 608 3696 1604
rect 3892 0 3960 312
rect 3892 608 3960 1604
rect 4156 0 4224 312
rect 4156 608 4224 1604
rect 4420 0 4488 312
rect 4420 608 4488 1604
rect 4684 0 4752 312
rect 4684 608 4752 1604
rect 4948 0 5016 312
rect 4948 608 5016 1604
rect 5212 0 5280 312
rect 5212 608 5280 1604
rect 5476 0 5544 312
rect 5476 608 5544 1604
rect 7852 0 7920 312
rect 7852 608 7920 1604
rect 8116 0 8184 312
rect 8116 608 8184 1604
rect 8380 0 8448 312
rect 8380 608 8448 1604
rect 8644 0 8712 312
rect 8644 608 8712 1604
rect 328 0 396 1536
rect 592 0 660 1536
rect 856 0 924 1536
rect 1120 0 1188 1536
rect 1384 0 1452 1536
rect 1648 0 1716 1536
rect 1912 0 1980 1536
rect 2176 0 2244 1536
rect 2440 0 2508 1536
rect 2704 0 2772 1536
rect 2968 0 3036 1536
rect 3232 0 3300 1536
rect 3496 0 3564 1536
rect 3760 0 3828 1536
rect 4024 0 4092 1536
rect 4288 0 4356 1536
rect 4552 0 4620 1536
rect 4816 0 4884 1536
rect 5080 0 5148 1536
rect 5344 0 5412 1536
rect 5608 0 5676 1536
rect 5872 0 5940 1536
rect 6136 0 6204 1536
rect 6400 0 6468 1536
rect 6664 0 6732 1536
rect 6928 0 6996 1536
rect 7192 0 7260 1536
rect 7456 0 7524 1536
rect 7720 0 7788 1536
rect 7984 0 8052 1536
rect 8248 0 8316 1536
rect 8512 0 8580 1536
rect 8908 0 8976 1604
rect 8776 0 8844 1604
rect 328 0 8908 68
rect 328 1536 8908 1604
<< m4 >>
rect 196 0 264 1604
rect 460 0 528 1604
rect 724 0 792 1604
rect 988 0 1056 1604
rect 1252 0 1320 1604
rect 1516 0 1584 1604
rect 1780 0 1848 1604
rect 2044 0 2112 1604
rect 2308 0 2376 1604
rect 2572 0 2640 1604
rect 2836 0 2904 1604
rect 3100 0 3168 1604
rect 3364 0 3432 1604
rect 3628 0 3696 1604
rect 3892 0 3960 1604
rect 4156 0 4224 1604
rect 4420 0 4488 1604
rect 4684 0 4752 1604
rect 4948 0 5016 1604
rect 5212 0 5280 1604
rect 5476 0 5544 1604
rect 5740 0 5808 1604
rect 6004 0 6072 1604
rect 6268 0 6336 1604
rect 6532 0 6600 1604
rect 6796 0 6864 1604
rect 7060 0 7128 1604
rect 7324 0 7392 1604
rect 7588 0 7656 1604
rect 7852 0 7920 1604
rect 8116 0 8184 1604
rect 8380 0 8448 1604
rect 8644 0 8712 1604
rect 8908 0 8976 1604
rect 196 0 8908 68
rect 196 1536 8908 1604
<< m3 >>
rect 328 0 396 1604
rect 460 132 528 1472
rect 592 0 660 1604
rect 724 132 792 1472
rect 856 0 924 1604
rect 988 132 1056 1472
rect 1120 0 1188 1604
rect 1252 132 1320 1472
rect 1384 0 1452 1604
rect 1516 132 1584 1472
rect 1648 0 1716 1604
rect 1780 132 1848 1472
rect 1912 0 1980 1604
rect 2044 132 2112 1472
rect 2176 0 2244 1604
rect 2308 132 2376 1472
rect 2440 0 2508 1604
rect 2572 132 2640 1472
rect 2704 0 2772 1604
rect 2836 132 2904 1472
rect 2968 0 3036 1604
rect 3100 132 3168 1472
rect 3232 0 3300 1604
rect 3364 132 3432 1472
rect 3496 0 3564 1604
rect 3628 132 3696 1472
rect 3760 0 3828 1604
rect 3892 132 3960 1472
rect 4024 0 4092 1604
rect 4156 132 4224 1472
rect 4288 0 4356 1604
rect 4420 132 4488 1472
rect 4552 0 4620 1604
rect 4684 132 4752 1472
rect 4816 0 4884 1604
rect 4948 132 5016 1472
rect 5080 0 5148 1604
rect 5212 132 5280 1472
rect 5344 0 5412 1604
rect 5476 132 5544 1472
rect 5608 0 5676 1604
rect 5740 132 5808 1472
rect 5872 0 5940 1604
rect 6004 132 6072 1472
rect 6136 0 6204 1604
rect 6268 132 6336 1472
rect 6400 0 6468 1604
rect 6532 132 6600 1472
rect 6664 0 6732 1604
rect 6796 132 6864 1472
rect 6928 0 6996 1604
rect 7060 132 7128 1472
rect 7192 0 7260 1604
rect 7324 132 7392 1472
rect 7456 0 7524 1604
rect 7588 132 7656 1472
rect 7720 0 7788 1604
rect 7852 132 7920 1472
rect 7984 0 8052 1604
rect 8116 132 8184 1472
rect 8248 0 8316 1604
rect 8380 132 8448 1472
rect 8512 0 8580 1604
rect 8644 132 8712 1472
rect 8908 0 8976 1604
rect 8776 0 8844 1604
rect 328 0 8776 68
rect 328 1536 8776 1604
<< m2 >>
rect 460 132 528 1472
rect 724 132 792 1472
rect 988 132 1056 1472
rect 1252 132 1320 1472
rect 1516 132 1584 1472
rect 1780 132 1848 1472
rect 2044 132 2112 1472
rect 2308 132 2376 1472
rect 2572 132 2640 1472
rect 2836 132 2904 1472
rect 3100 132 3168 1472
rect 3364 132 3432 1472
rect 3628 132 3696 1472
rect 3892 132 3960 1472
rect 4156 132 4224 1472
rect 4420 132 4488 1472
rect 4684 132 4752 1472
rect 4948 132 5016 1472
rect 5212 132 5280 1472
rect 5476 132 5544 1472
rect 5740 132 5808 1472
rect 6004 132 6072 1472
rect 6268 132 6336 1472
rect 6532 132 6600 1472
rect 6796 132 6864 1472
rect 7060 132 7128 1472
rect 7324 132 7392 1472
rect 7588 132 7656 1472
rect 7852 132 7920 1472
rect 8116 132 8184 1472
rect 8380 132 8448 1472
rect 8644 132 8712 1472
rect 8908 0 8976 1604
<< locali >>
rect 0 426 8776 494
rect 0 198 8776 266
rect 0 1338 8776 1406
rect 0 654 8776 722
rect 0 1110 8776 1178
rect 0 882 8776 950
use RM1 XRES1A
transform 1 0 200 0 1 198
box 200 198 320 198
use RM1 XRES1B
transform 1 0 200 0 1 1338
box 200 1338 320 1338
use RM1 XRES2
transform 1 0 200 0 1 654
box 200 654 320 654
use RM1 XRES4
transform 1 0 200 0 1 1110
box 200 1110 320 1110
use RM1 XRES8
transform 1 0 200 0 1 882
box 200 882 320 882
use RM1 XRES16
transform 1 0 200 0 1 426
box 200 426 320 426
use cut_M2M5_1x2 
transform 1 0 8908 0 1 602
box 8908 602 8976 802
use cut_M1M4_1x2 
transform 1 0 2308 0 1 132
box 2308 132 2376 332
use cut_M1M4_1x2 
transform 1 0 6796 0 1 1272
box 6796 1272 6864 1472
use cut_M1M4_1x2 
transform 1 0 2572 0 1 588
box 2572 588 2640 788
use cut_M1M4_1x2 
transform 1 0 6532 0 1 588
box 6532 588 6600 788
use cut_M1M4_1x2 
transform 1 0 2044 0 1 1044
box 2044 1044 2112 1244
use cut_M1M4_1x2 
transform 1 0 2836 0 1 1044
box 2836 1044 2904 1244
use cut_M1M4_1x2 
transform 1 0 6268 0 1 1044
box 6268 1044 6336 1244
use cut_M1M4_1x2 
transform 1 0 7060 0 1 1044
box 7060 1044 7128 1244
use cut_M1M4_1x2 
transform 1 0 1516 0 1 816
box 1516 816 1584 1016
use cut_M1M4_1x2 
transform 1 0 1780 0 1 816
box 1780 816 1848 1016
use cut_M1M4_1x2 
transform 1 0 3100 0 1 816
box 3100 816 3168 1016
use cut_M1M4_1x2 
transform 1 0 3364 0 1 816
box 3364 816 3432 1016
use cut_M1M4_1x2 
transform 1 0 5740 0 1 816
box 5740 816 5808 1016
use cut_M1M4_1x2 
transform 1 0 6004 0 1 816
box 6004 816 6072 1016
use cut_M1M4_1x2 
transform 1 0 7324 0 1 816
box 7324 816 7392 1016
use cut_M1M4_1x2 
transform 1 0 7588 0 1 816
box 7588 816 7656 1016
use cut_M1M4_1x2 
transform 1 0 460 0 1 360
box 460 360 528 560
use cut_M1M4_1x2 
transform 1 0 724 0 1 360
box 724 360 792 560
use cut_M1M4_1x2 
transform 1 0 988 0 1 360
box 988 360 1056 560
use cut_M1M4_1x2 
transform 1 0 1252 0 1 360
box 1252 360 1320 560
use cut_M1M4_1x2 
transform 1 0 3628 0 1 360
box 3628 360 3696 560
use cut_M1M4_1x2 
transform 1 0 3892 0 1 360
box 3892 360 3960 560
use cut_M1M4_1x2 
transform 1 0 4156 0 1 360
box 4156 360 4224 560
use cut_M1M4_1x2 
transform 1 0 4420 0 1 360
box 4420 360 4488 560
use cut_M1M4_1x2 
transform 1 0 4684 0 1 360
box 4684 360 4752 560
use cut_M1M4_1x2 
transform 1 0 4948 0 1 360
box 4948 360 5016 560
use cut_M1M4_1x2 
transform 1 0 5212 0 1 360
box 5212 360 5280 560
use cut_M1M4_1x2 
transform 1 0 5476 0 1 360
box 5476 360 5544 560
use cut_M1M4_1x2 
transform 1 0 7852 0 1 360
box 7852 360 7920 560
use cut_M1M4_1x2 
transform 1 0 8116 0 1 360
box 8116 360 8184 560
use cut_M1M4_1x2 
transform 1 0 8380 0 1 360
box 8380 360 8448 560
use cut_M1M4_1x2 
transform 1 0 8644 0 1 360
box 8644 360 8712 560
<< labels >>
flabel m3 s 328 0 396 1604 0 FreeSans 400 0 0 0 CTOP
port 1 nsew
flabel m1 s 328 0 8908 68 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 0 198 200 266 0 FreeSans 400 0 0 0 C1A
port 3 nsew
flabel locali s 0 1338 200 1406 0 FreeSans 400 0 0 0 C1B
port 4 nsew
flabel locali s 0 654 200 722 0 FreeSans 400 0 0 0 C2
port 5 nsew
flabel locali s 0 1110 200 1178 0 FreeSans 400 0 0 0 C4
port 6 nsew
flabel locali s 0 882 200 950 0 FreeSans 400 0 0 0 C8
port 7 nsew
flabel locali s 0 426 200 494 0 FreeSans 400 0 0 0 C16
port 8 nsew
<< end >>
