magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 4056 5760
<< locali >>
rect 3432 384 3672 5376
rect 384 384 3672 624
rect 384 5136 3672 5376
rect 384 384 624 5376
rect 3432 384 3672 5376
rect 3816 0 4056 5760
rect 0 0 4056 240
rect 0 5520 4056 5760
rect 0 0 240 5760
rect 3816 0 4056 5760
rect 1200 2322 1368 2382
rect 1368 1530 1632 1590
rect 1200 3026 1368 3086
rect 1368 1530 1428 3086
<< m1 >>
rect 1200 2674 1368 2734
rect 1368 2410 1632 2470
rect 1368 2410 1428 2734
rect 1200 3378 1368 3438
rect 1368 3994 1632 4054
rect 1200 4786 1368 4846
rect 1368 3378 1428 4846
rect 972 1266 1200 1326
rect 972 3230 1584 3290
rect 972 3670 1152 3730
rect 972 1266 1032 3730
rect 1524 3290 1632 3350
rect 1092 3730 1200 3790
<< m3 >>
rect 1516 384 1732 4992
rect 2308 768 2524 5760
<< m2 >>
rect 3840 2762 4056 2822
rect 0 1618 216 1678
rect 3840 4874 4056 4934
rect 0 4082 216 4142
rect 0 1618 216 1678
rect 952 1618 1200 1694
rect 108 1618 952 1694
rect 952 1618 1028 1694
rect 0 4082 216 4142
rect 952 4082 1200 4158
rect 108 4082 952 4158
rect 952 4082 1028 4158
rect 3840 2762 4056 2822
rect 1632 2762 1804 2838
rect 1804 2762 3948 2838
rect 1804 2762 1880 2838
rect 3840 4874 4056 4934
rect 1632 4874 1804 4950
rect 1804 4874 3948 4950
rect 1804 4874 1880 4950
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV xa00
transform 1 0 768 0 1 768
box 768 768 3288 1120
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV xa10
transform 1 0 768 0 1 1120
box 768 1120 3288 2176
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa20
transform 1 0 768 0 1 2176
box 768 2176 3288 2528
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa2a0
transform 1 0 768 0 1 2528
box 768 2528 3288 2880
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NRX1_CV xa30
transform 1 0 768 0 1 2880
box 768 2880 3288 3584
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV xa50
transform 1 0 768 0 1 3584
box 768 3584 3288 4640
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa60
transform 1 0 768 0 1 4640
box 768 4640 3288 4992
use cut_M1M2_2x1 
transform 1 0 1092 0 1 2674
box 1092 2674 1276 2742
use cut_M1M2_2x1 
transform 1 0 1524 0 1 2410
box 1524 2410 1708 2478
use cut_M1M2_2x1 
transform 1 0 1092 0 1 3378
box 1092 3378 1276 3446
use cut_M1M2_2x1 
transform 1 0 1524 0 1 3994
box 1524 3994 1708 4062
use cut_M1M2_2x1 
transform 1 0 1092 0 1 4786
box 1092 4786 1276 4854
use cut_M1M2_2x1 
transform 1 0 1124 0 1 1266
box 1124 1266 1308 1334
use cut_M1M2_2x1 
transform 1 0 1556 0 1 3290
box 1556 3290 1740 3358
use cut_M1M2_2x1 
transform 1 0 1124 0 1 3730
box 1124 3730 1308 3798
use cut_M1M4_2x1 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 
transform 1 0 2316 0 1 5520
box 2316 5520 2516 5596
use cut_M1M3_2x1 
transform 1 0 1108 0 1 1618
box 1108 1618 1308 1694
use cut_M1M3_2x1 
transform 1 0 1108 0 1 4082
box 1108 4082 1308 4158
use cut_M1M3_2x1 
transform 1 0 1524 0 1 2762
box 1524 2762 1724 2838
use cut_M1M3_2x1 
transform 1 0 1524 0 1 4874
box 1524 4874 1724 4950
<< labels >>
flabel locali s 3432 384 3672 5376 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 3816 0 4056 5760 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 3840 2762 4056 2822 0 FreeSans 400 0 0 0 CP_UP_N
port 2 nsew
flabel m2 s 0 1618 216 1678 0 FreeSans 400 0 0 0 CK_REF
port 3 nsew
flabel m2 s 3840 4874 4056 4934 0 FreeSans 400 0 0 0 CP_DOWN
port 4 nsew
flabel m2 s 0 4082 216 4142 0 FreeSans 400 0 0 0 CK_FB
port 5 nsew
<< end >>
