magic
tech sky130A
magscale 1 2
timestamp 1660661870
<< checkpaint >>
rect 0 0 200 76
<< m3 >>
rect 0 0 200 76
<< v3 >>
rect 12 6 76 70
rect 124 6 188 70
<< m4 >>
rect 0 0 200 76
<< labels >>
<< end >>
