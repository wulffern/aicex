
.subckt NCHDLCM D G S B
M0 N0 G  S B NCHDL2
M1 N1 G  N0 B NCHDL2
M2 N2 G  N1 B NCHDL2
M3 N3 G  N2 B NCHDL2
M4 N4 G  N3 B NCHDL2
M5 N5 G  N4 B NCHDL2
M6 N6 G  N5 B NCHDL2
M7 N7 G  N6 B NCHDL2
M8 D G N7  B NCHDL2
.ends

.subckt PCHDLCM D G S B
M0 N0 G  S B PCHDL2
M7 D G N0  B PCHDL2
.ends


.subckt NCHDLA D G S B
M0 D G  S B NCHDL2
M1 S G  D B NCHDL2
.ends

.subckt PCHDLA D G S B
M0 D G S B PCHDL2
M1 S G D B PCHDL2
M2 D G S B PCHDL2
M3 S G D B PCHDL2
M4 D G S B PCHDL2
M5 S G D B PCHDL2
M6 D G S B PCHDL2
M7 S G D B PCHDL2
.ends

.subckt NCHDLCM2 D G S B
M0 D G  S B NCHDLCM
M1 S G  D B NCHDLCM
.ends

.subckt PCHDLCM2 D G S B
M0 D G  S B PCHDLCM
M1 S G D B PCHDLCM
.ends

.subckt PCHDLCM2 D G S B
M0 D G  S B PCHDLCM
M1 S G D B PCHDLCM
.ends

.subckt CPCHDLCM2 D G CG S CS B
M0 CS G S B PCHDLCM2
M1 D CG CS B PCHDLA
.ends

.subckt CNCHDLCM2 D G CG S CS B
M0 CS G S B NCHDLCM2
M1 D CG CS B NCHDLA
.ends
