magic
tech sky130A
magscale 1 2
timestamp 1661983200
<< checkpaint >>
rect 0 0 3888 2860
<< locali >>
rect 3384 2750 3960 2970
rect -72 2750 504 2970
use SUNTR_RES8 XA1
transform 1 0 0 0 1 0
box 0 0 3888 2860
<< labels >>
flabel locali s 3384 2750 3960 2970 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s -72 2750 504 2970 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
