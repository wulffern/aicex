magic
tech sky130A
magscale 1 2
timestamp 1661001370
<< checkpaint >>
rect -768 -768 13368 6252
<< locali >>
rect 12744 -384 12984 5664
rect -384 -384 12984 -144
rect -384 5424 12984 5664
rect -384 -384 -144 5664
rect 12744 -384 12984 5664
rect 13128 -768 13368 6048
rect -768 -768 13368 -528
rect -768 5808 13368 6048
rect -768 -768 -528 6048
rect 13128 -768 13368 6048
rect -768 6192 13368 6252
rect -768 6192 13368 6252
rect 756 5162 972 5222
rect 10404 498 10620 558
<< m3 >>
rect 748 -384 964 5280
rect 4076 -384 4292 5280
rect 5788 -384 6004 5280
rect 9116 -384 9332 5280
rect 10828 -384 11044 5280
rect 1540 -768 1756 5280
rect 3284 -768 3500 5280
rect 6580 -768 6796 5280
rect 8324 -768 8540 5280
rect 11620 -768 11836 5280
rect 394 4018 470 6252
rect 4570 4018 4646 6252
rect 5434 4018 5510 6252
rect 9610 4018 9686 6252
rect 10474 4018 10550 6252
<< m1 >>
rect 864 4810 1032 4870
rect 1032 1614 2040 1674
rect 1032 1554 1092 4870
rect 1980 1554 2088 1614
rect 5904 4810 6072 4870
rect 6072 1614 7080 1674
rect 6072 1554 6132 4870
rect 7020 1554 7128 1614
rect 10944 4810 11112 4870
rect 11112 1614 12120 1674
rect 11112 1554 11172 4870
rect 12060 1554 12168 1614
rect 3948 4810 4176 4870
rect 3000 1614 3948 1674
rect 3948 1554 4008 4870
rect 2952 1554 3060 1614
rect 8988 4810 9216 4870
rect 8040 1614 8988 1674
rect 8988 1554 9048 4870
rect 7992 1554 8100 1614
<< m2 >>
rect 4608 498 4988 574
rect 4988 5238 5856 5314
rect 4988 498 5064 5314
rect 5796 5162 5904 5238
rect 9648 498 10028 574
rect 10028 5238 10896 5314
rect 10028 498 10104 5314
rect 10836 5162 10944 5238
rect 480 574 2468 650
rect 2468 5238 4128 5314
rect 2468 498 2544 5314
rect 432 498 540 574
rect 4068 5162 4176 5238
rect 5520 574 7508 650
rect 7508 5238 9168 5314
rect 7508 498 7584 5314
rect 5472 498 5580 574
rect 9108 5162 9216 5238
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xc0
transform 1 0 0 0 1 0
box 0 0 2520 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xd0
transform -1 0 5040 0 1 0
box 5040 0 7560 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xe0
transform 1 0 5040 0 1 0
box 5040 0 7560 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xf0
transform -1 0 10080 0 1 0
box 10080 0 12600 5280
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xg0
transform 1 0 10080 0 1 0
box 10080 0 12600 5280
use cut_M1M4_2x1 
transform 1 0 756 0 1 -384
box 756 -384 956 -308
use cut_M1M4_2x1 
transform 1 0 4084 0 1 -384
box 4084 -384 4284 -308
use cut_M1M4_2x1 
transform 1 0 5796 0 1 -384
box 5796 -384 5996 -308
use cut_M1M4_2x1 
transform 1 0 9124 0 1 -384
box 9124 -384 9324 -308
use cut_M1M4_2x1 
transform 1 0 10836 0 1 -384
box 10836 -384 11036 -308
use cut_M1M4_2x1 
transform 1 0 1548 0 1 -768
box 1548 -768 1748 -692
use cut_M1M4_2x1 
transform 1 0 3292 0 1 -768
box 3292 -768 3492 -692
use cut_M1M4_2x1 
transform 1 0 6588 0 1 -768
box 6588 -768 6788 -692
use cut_M1M4_2x1 
transform 1 0 8332 0 1 -768
box 8332 -768 8532 -692
use cut_M1M4_2x1 
transform 1 0 11628 0 1 -768
box 11628 -768 11828 -692
use cut_M2M4_2x1 
transform 1 0 332 0 1 4018
box 332 4018 532 4094
use cut_M1M4_2x1 
transform 1 0 332 0 1 6192
box 332 6192 532 6268
use cut_M2M4_2x1 
transform 1 0 4508 0 1 4018
box 4508 4018 4708 4094
use cut_M1M4_2x1 
transform 1 0 4508 0 1 6192
box 4508 6192 4708 6268
use cut_M2M4_2x1 
transform 1 0 5372 0 1 4018
box 5372 4018 5572 4094
use cut_M1M4_2x1 
transform 1 0 5372 0 1 6192
box 5372 6192 5572 6268
use cut_M2M4_2x1 
transform 1 0 9548 0 1 4018
box 9548 4018 9748 4094
use cut_M1M4_2x1 
transform 1 0 9548 0 1 6192
box 9548 6192 9748 6268
use cut_M2M4_2x1 
transform 1 0 10412 0 1 4018
box 10412 4018 10612 4094
use cut_M1M4_2x1 
transform 1 0 10412 0 1 6192
box 10412 6192 10612 6268
use cut_M1M2_2x1 
transform 1 0 1980 0 1 1554
box 1980 1554 2164 1622
use cut_M1M2_2x1 
transform 1 0 7020 0 1 1554
box 7020 1554 7204 1622
use cut_M1M2_2x1 
transform 1 0 12060 0 1 1554
box 12060 1554 12244 1622
use cut_M1M2_2x1 
transform 1 0 2876 0 1 1554
box 2876 1554 3060 1622
use cut_M1M2_2x1 
transform 1 0 7916 0 1 1554
box 7916 1554 8100 1622
use cut_M1M3_2x1 
transform 1 0 4500 0 1 498
box 4500 498 4700 574
use cut_M1M3_2x1 
transform 1 0 5796 0 1 5162
box 5796 5162 5996 5238
use cut_M1M3_2x1 
transform 1 0 9540 0 1 498
box 9540 498 9740 574
use cut_M1M3_2x1 
transform 1 0 10836 0 1 5162
box 10836 5162 11036 5238
use cut_M1M3_2x1 
transform 1 0 324 0 1 498
box 324 498 524 574
use cut_M1M3_2x1 
transform 1 0 4068 0 1 5162
box 4068 5162 4268 5238
use cut_M1M3_2x1 
transform 1 0 5364 0 1 498
box 5364 498 5564 574
use cut_M1M3_2x1 
transform 1 0 9108 0 1 5162
box 9108 5162 9308 5238
<< labels >>
flabel locali s 12744 -384 12984 5664 0 FreeSans 400 0 0 0 AVSS
port 5 nsew
flabel locali s 13128 -768 13368 6048 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s -768 6192 13368 6252 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew
flabel locali s 756 5162 972 5222 0 FreeSans 400 0 0 0 CK_FB
port 2 nsew
flabel locali s 10404 498 10620 558 0 FreeSans 400 0 0 0 CK
port 3 nsew
<< end >>
