magic
tech sky130A
magscale 1 2
timestamp 1658600916
<< checkpaint >>
rect 0 0 152 0
<< m3 >>
rect 0 0 76 76
rect 0 0 76 76
rect 76 0 228 76
rect 76 0 228 76
<< rm3 >>
rect 76 0 152 76
<< labels >>
flabel m3 s 0 0 76 76 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel m3 s 76 0 228 76 0 FreeSans 400 0 0 0 B
port 2 nsew
<< end >>
