magic
tech sky130A
magscale 1 2
timestamp 1660117866
<< checkpaint >>
rect -768 -768 13944 11328
<< locali >>
rect 13320 -384 13560 10944
rect -384 -384 13560 -144
rect -384 10704 13560 10944
rect -384 -384 -144 10944
rect 13320 -384 13560 10944
rect 756 -384 972 118
rect -108 -384 108 220
rect 756 -384 972 118
rect -108 -384 108 220
rect -108 -384 108 1980
rect -108 -384 108 2508
rect 13704 -768 13944 11328
rect -768 -768 13944 -528
rect -768 11088 13944 11328
rect -768 -768 -528 11328
rect 13704 -768 13944 11328
rect 2376 -768 2592 118
rect 1512 -768 1728 220
rect 2376 -768 2592 118
rect 1512 -768 1728 220
rect 864 1642 1032 1702
rect 864 1818 1032 1878
rect 864 2346 1032 2406
rect 1032 1642 1092 2406
rect 2484 58 2652 118
rect 2484 1290 2652 1350
rect 2484 2522 2652 2582
rect 2484 3754 2652 3814
rect 2484 4986 2652 5046
rect 2484 6218 2652 6278
rect 2484 7450 2652 7510
rect 2484 8682 2652 8742
rect 2652 58 2712 8742
rect 324 146 540 206
rect 324 2434 540 2494
rect 2376 2698 2592 2758
rect 324 1906 540 1966
<< m3 >>
rect 8028 -384 8244 44
rect 2484 2698 2664 2774
rect 2484 3930 2664 4006
rect 2484 5162 2664 5238
rect 2484 6394 2664 6470
rect 2484 7626 2664 7702
rect 2484 8858 2664 8934
rect 2664 836 8136 912
rect 2664 1892 8136 1968
rect 2664 2948 8136 3024
rect 2664 4004 8136 4080
rect 2664 5060 8136 5136
rect 2664 6116 8136 6192
rect 2664 7172 8136 7248
rect 2664 8228 8136 8304
rect 2664 9284 8136 9360
rect 2664 10340 8136 10416
rect 2664 836 2740 10416
rect 8136 -44 13428 32
rect 8136 1012 13428 1088
rect 8136 2068 13428 2144
rect 8136 3124 13428 3200
rect 8136 4180 13428 4256
rect 8136 5236 13428 5312
rect 8136 6292 13428 6368
rect 8136 7348 13428 7424
rect 8136 8404 13428 8480
rect 8136 9460 13428 9536
rect 13428 -44 13504 9536
<< m1 >>
rect 2052 8770 2220 8830
rect 2220 234 2484 294
rect 2052 2610 2220 2670
rect 2052 3842 2220 3902
rect 2052 5074 2220 5134
rect 2052 6306 2220 6366
rect 2052 7538 2220 7598
rect 864 2522 2220 2582
rect 2220 234 2280 8838
<< m2 >>
rect 2052 146 2224 222
rect 864 1994 2224 2070
rect 2224 1466 2484 1542
rect 2052 1378 2224 1454
rect 2224 146 2300 2070
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa1
transform 1 0 0 0 1 0
box 0 0 1260 1760
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa2
transform 1 0 0 0 1 1760
box 0 1760 1260 2288
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa4
transform 1 0 0 0 1 2288
box 0 2288 1260 2816
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc1
transform -1 0 2880 0 1 0
box 2880 0 4140 1232
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc2
transform -1 0 2880 0 1 1232
box 2880 1232 4140 2464
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_0
transform -1 0 2880 0 1 2464
box 2880 2464 4140 3696
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_1
transform -1 0 2880 0 1 3696
box 2880 3696 4140 4928
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_2
transform -1 0 2880 0 1 4928
box 2880 4928 4140 6160
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_3
transform -1 0 2880 0 1 6160
box 2880 6160 4140 7392
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_4
transform -1 0 2880 0 1 7392
box 2880 7392 4140 8624
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_5
transform -1 0 2880 0 1 8624
box 2880 8624 4140 9856
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd20
transform 1 0 3024 0 1 0
box 3024 0 13176 1056
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd30
transform 1 0 3024 0 1 1056
box 3024 1056 13176 2112
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd31
transform 1 0 3024 0 1 2112
box 3024 2112 13176 3168
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd32
transform 1 0 3024 0 1 3168
box 3024 3168 13176 4224
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd33
transform 1 0 3024 0 1 4224
box 3024 4224 13176 5280
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd34
transform 1 0 3024 0 1 5280
box 3024 5280 13176 6336
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd35
transform 1 0 3024 0 1 6336
box 3024 6336 13176 7392
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd36
transform 1 0 3024 0 1 7392
box 3024 7392 13176 8448
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd37
transform 1 0 3024 0 1 8448
box 3024 8448 13176 9504
use ../../sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd38
transform 1 0 3024 0 1 9504
box 3024 9504 13176 10560
use cut_M1M4_2x1 
transform 1 0 8036 0 1 -384
box 8036 -384 8236 -308
use cut_M1M2_2x1 
transform 1 0 1944 0 1 8770
box 1944 8770 2128 8838
use cut_M1M2_2x1 
transform 1 0 2376 0 1 234
box 2376 234 2560 302
use cut_M1M2_2x1 
transform 1 0 1944 0 1 2610
box 1944 2610 2128 2678
use cut_M1M2_2x1 
transform 1 0 1944 0 1 3842
box 1944 3842 2128 3910
use cut_M1M2_2x1 
transform 1 0 1944 0 1 5074
box 1944 5074 2128 5142
use cut_M1M2_2x1 
transform 1 0 1944 0 1 6306
box 1944 6306 2128 6374
use cut_M1M2_2x1 
transform 1 0 1944 0 1 7538
box 1944 7538 2128 7606
use cut_M1M2_2x1 
transform 1 0 756 0 1 2522
box 756 2522 940 2590
use cut_M1M3_2x1 
transform 1 0 1944 0 1 146
box 1944 146 2144 222
use cut_M1M3_2x1 
transform 1 0 756 0 1 1994
box 756 1994 956 2070
use cut_M1M3_2x1 
transform 1 0 2376 0 1 1466
box 2376 1466 2576 1542
use cut_M1M3_2x1 
transform 1 0 1944 0 1 1378
box 1944 1378 2144 1454
use cut_M1M3_2x1 
transform 1 0 2376 0 1 1466
box 2376 1466 2576 1542
use cut_M1M3_2x1 
transform 1 0 1944 0 1 1378
box 1944 1378 2144 1454
use cut_M1M4_2x1 
transform 1 0 2376 0 1 2698
box 2376 2698 2576 2774
use cut_M1M4_2x1 
transform 1 0 2376 0 1 3930
box 2376 3930 2576 4006
use cut_M1M4_2x1 
transform 1 0 2376 0 1 5162
box 2376 5162 2576 5238
use cut_M1M4_2x1 
transform 1 0 2376 0 1 6394
box 2376 6394 2576 6470
use cut_M1M4_2x1 
transform 1 0 2376 0 1 7626
box 2376 7626 2576 7702
use cut_M1M4_2x1 
transform 1 0 2376 0 1 8858
box 2376 8858 2576 8934
<< labels >>
flabel locali s 13320 -384 13560 10944 0 FreeSans 400 0 0 0 AVSS
port 3 nsew
flabel locali s 13704 -768 13944 11328 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 VBN
port 2 nsew
flabel locali s 324 2434 540 2494 0 FreeSans 400 0 0 0 VI
port 4 nsew
flabel locali s 2376 2698 2592 2758 0 FreeSans 400 0 0 0 VO
port 5 nsew
flabel locali s 324 1906 540 1966 0 FreeSans 400 0 0 0 VFB
port 6 nsew
<< end >>
