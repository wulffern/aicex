magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 3840
<< locali >>
rect 1740 450 1894 510
rect 1740 2690 1894 2750
rect 1740 3650 1894 3710
rect 1894 450 1954 3710
rect 390 1670 514 1730
rect 514 1490 720 1550
rect 514 1490 574 1730
rect 390 1730 450 1790
rect 360 3330 514 3390
rect 514 1810 720 1870
rect 514 1810 574 3390
rect 360 2370 514 2430
rect 514 1810 720 1870
rect 514 1810 574 2430
rect 146 770 360 830
rect 146 3010 360 3070
rect 146 770 206 3070
rect 270 2050 450 2110
rect 1650 3650 1830 3710
rect 270 450 450 510
rect 270 3010 450 3070
rect 630 2770 810 2830
rect 630 3730 810 3790
rect 1290 690 1470 750
<< m1 >>
rect 360 1090 514 1150
rect 360 2050 514 2110
rect 514 1090 574 2118
rect 146 450 360 510
rect 146 3650 360 3710
rect 146 2690 360 2750
rect 146 450 206 3718
<< m3 >>
rect 1290 0 1474 3840
rect 630 0 814 3840
rect 1290 0 1474 3840
rect 630 0 814 3840
use TAPCELLB_CV XA0
transform 1 0 0 0 1 0
box 0 0 2100 320
use SAREMX1_CV XA1
transform 1 0 0 0 1 320
box 0 320 2100 1600
use IVX1_CV XA2
transform 1 0 0 0 1 1600
box 0 1600 2100 1920
use SARLTX1_CV XA4
transform 1 0 0 0 1 1920
box 0 1920 2100 2880
use SARLTX1_CV XA5
transform 1 0 0 0 1 2880
box 0 2880 2100 3840
use cut_M1M2_2x1 
transform 1 0 266 0 1 1090
box 266 1090 450 1158
use cut_M1M2_2x1 
transform 1 0 266 0 1 2050
box 266 2050 450 2118
use cut_M1M2_2x1 
transform 1 0 270 0 1 450
box 270 450 454 518
use cut_M1M2_2x1 
transform 1 0 270 0 1 3650
box 270 3650 454 3718
use cut_M1M2_2x1 
transform 1 0 270 0 1 2690
box 270 2690 454 2758
<< labels >>
flabel locali s 270 2050 450 2110 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1650 3650 1830 3710 0 FreeSans 400 0 0 0 RST_N
port 2 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 270 3010 450 3070 0 FreeSans 400 0 0 0 CMP_ON
port 4 nsew
flabel locali s 630 2770 810 2830 0 FreeSans 400 0 0 0 CHL_OP
port 5 nsew
flabel locali s 630 3730 810 3790 0 FreeSans 400 0 0 0 CHL_ON
port 6 nsew
flabel locali s 1290 690 1470 750 0 FreeSans 400 0 0 0 ENO
port 7 nsew
flabel m3 s 1290 0 1474 3840 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 3840 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
