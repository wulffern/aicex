*RPLY_BIAS_SKY130A/RPLY_BIAS
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_BIAS_lpe.spi
#else
.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_10_lpe.spi
*.include ../../../../sun_tr_sky130nm/work/lpe/SUNTR_CAP_20_lpe.spi
.include ../../../work/xsch/RPLY_BIAS.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12 method=gear
#else
.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15 method=gear
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param T_END = {10u}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VPWR  PWRUP_1V8  VSS  pwl 0 0 20n 0 20.1n {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------

XDUT VDD_1V8 VSS PWRUP_1V8 LPO LPO IBP_1U<3>,IBP_1U<2>,IBP_1U<1>,IBP_1U<0> RPLY_BIAS
*-----------------------------------------------------------------
* STASH
*-----------------------------------------------------------------

V3 IBP_1U<3> 0 dc {AVDD/2}
V2 IBP_1U<2> 0 dc {AVDD/2}
V1 IBP_1U<1> 0 dc {AVDD/2}
V0 IBP_1U<0> 0 dc {AVDD/2}

B1 D_VD 0 v=v(XDUT.VR1)-v(XDUT.VD2)

B4 V_OFF 0 v=v(XDUT.VR1)-v(XDUT.VD1)

B2 D_VD_REF 0 v=1.38062e-23/1.60219e-19*(temper + 273.15)*ln(64)
B3 D_VD_ERR 0 v=v(D_VD)-v(D_VD_REF)
*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------
.measure tran ibp_1u FIND i(V1) AT={T_END}
.measure tran ivdd FIND i(VDD) AT={T_END}
.measure tran vd1 FIND v(XDUT.VD1) AT={T_END}
.measure tran vd2 FIND v(XDUT.VD2) AT={T_END}
.measure tran vr1 FIND v(XDUT.VR1) AT={T_END}
.measure tran m_offset FIND v(V_OFF) AT={T_END}
.measure tran dvd FIND v(D_VD) AT={T_END}
.measure tran dvdref FIND v(D_VD_REF) AT={T_END}
.measure tran dvderr FIND v(D_VD_ERR) AT={T_END}

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.probe v(VDD_1V8) v(VSS) v(PWRUP_1V8) v(LPI) v(LPO) v(IBP_1U) i(v1)
+ v(XDUT.VD1) v(XDUT.VD2) v(XDUT.VR1) v(D_VD) v(D_VD_REF) v(D_VD_ERR)
+ v(V_OFF) i(VDD)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

tran 10n 10.1u 1n
write
#ifdef Debug


*quit
#else

quit
#endif
.endc
