** sch_path:
*+ /Users/wulff/pro/aicex/ip/sun_pll_sky130nm/work/../design/SUN_PLL_SKY130NM/SUN_PLL_LPF.sch
.subckt SUN_PLL_LPF VLPF AVSS
*.ipin VLPF
*.ipin AVSS
xa3 VN1 VLPF AVSS SUNTR_RPPO_12k xoffset=0 yoffset=5 angle=0 M=1
xb1 VLPF AVSS CAP_LPF xoffset=0 yoffset=0 angle=0 M=1
xb2 VLPF AVSS CAP_LPF xoffset=0 yoffset=0 angle=0 M=1
xb3 VN1 AVSS CAP_LPF xoffset=0 yoffset=0 angle=0 M=5
.ends

* expanding   symbol:  SUN_PLL_SKY130NM/CAP_LPF.sym # of pins=2
** sym_path:
*+ /Users/wulff/Documents/pro/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/CAP_LPF.sym
** sch_path:
*+ /Users/wulff/Documents/pro/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/CAP_LPF.sch
.subckt CAP_LPF  A B   xoffset=0 yoffset=0 angle=0 M=1
*.iopin A
*.iopin B
R1 A NC0 sky130_fd_pr__res_generic_m1 W=0.4 L=0.4 m=1
R2 B NC1 sky130_fd_pr__res_generic_m1 W=0.4 L=0.4 m=1
.ends

.end
