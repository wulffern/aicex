* NGSPICE file created from SAR9B_CV.ext - technology: sky130A

.subckt SAR9B_CV SAR_IP SAR_IN SARN SARP DONE D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1>
+ D<0> EN CK_SAMPLE CK_SAMPLE_BSSW VREF AVDD AVSS
R0 XA0/CP0 XDAC1/XC128b<2>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R1 XA0/CP0 XDAC1/XC128b<2>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R2 XA0/CP0 XDAC1/XC128b<2>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R3 XA0/CP0 XDAC1/XC128b<2>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R4 XA0/CP0 XDAC1/XC128b<2>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R5 XA0/CP0 XDAC1/XC128b<2>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R6 XA2/CP0 XDAC1/X16ab/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R7 D<5> XDAC1/X16ab/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R8 D<5> XDAC1/X16ab/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R9 D<5> XDAC1/X16ab/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R10 D<5> XDAC1/X16ab/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R11 XA3/CP0 XDAC1/X16ab/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R12 XA1/CP0 XDAC1/XC64a<0>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R13 XA1/CP0 XDAC1/XC64a<0>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R14 XA1/CP0 XDAC1/XC64a<0>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R15 XA1/CP0 XDAC1/XC64a<0>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R16 XA1/CP0 XDAC1/XC64a<0>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R17 XA1/CP0 XDAC1/XC64a<0>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R18 XA0/CP1 XDAC1/XC0/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R19 XA0/CP1 XDAC1/XC0/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R20 XA0/CP1 XDAC1/XC0/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R21 XA0/CP1 XDAC1/XC0/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R22 XA0/CP1 XDAC1/XC0/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R23 XA0/CP1 XDAC1/XC0/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R24 XA0/CP0 XDAC1/XC1/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R25 XA0/CP0 XDAC1/XC1/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R26 XA0/CP0 XDAC1/XC1/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R27 XA0/CP0 XDAC1/XC1/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R28 XA0/CP0 XDAC1/XC1/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R29 XA0/CP0 XDAC1/XC1/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R30 D<7> XDAC1/XC64b<1>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R31 D<7> XDAC1/XC64b<1>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R32 D<7> XDAC1/XC64b<1>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R33 D<7> XDAC1/XC64b<1>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R34 D<7> XDAC1/XC64b<1>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R35 D<7> XDAC1/XC64b<1>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R36 XA0/CP1 XDAC1/XC128a<1>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R37 XA0/CP1 XDAC1/XC128a<1>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R38 XA0/CP1 XDAC1/XC128a<1>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R39 XA0/CP1 XDAC1/XC128a<1>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R40 XA0/CP1 XDAC1/XC128a<1>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R41 XA0/CP1 XDAC1/XC128a<1>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R42 D<6> XDAC1/XC32a<0>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R43 XDAC1/XC32a<0>/C1A AVSS sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R44 D<2> XDAC1/XC32a<0>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R45 D<1> XDAC1/XC32a<0>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R46 D<3> XDAC1/XC32a<0>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R47 D<4> XDAC1/XC32a<0>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R48 XA0/CN0 XDAC2/XC128b<2>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R49 XA0/CN0 XDAC2/XC128b<2>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R50 XA0/CN0 XDAC2/XC128b<2>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R51 XA0/CN0 XDAC2/XC128b<2>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R52 XA0/CN0 XDAC2/XC128b<2>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R53 XA0/CN0 XDAC2/XC128b<2>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R54 XA2/CN0 XDAC2/X16ab/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R55 XA3/CN1 XDAC2/X16ab/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R56 XA3/CN1 XDAC2/X16ab/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R57 XA3/CN1 XDAC2/X16ab/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R58 XA3/CN1 XDAC2/X16ab/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R59 XA3/CN0 XDAC2/X16ab/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R60 XA1/CN0 XDAC2/XC64a<0>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R61 XA1/CN0 XDAC2/XC64a<0>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R62 XA1/CN0 XDAC2/XC64a<0>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R63 XA1/CN0 XDAC2/XC64a<0>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R64 XA1/CN0 XDAC2/XC64a<0>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R65 XA1/CN0 XDAC2/XC64a<0>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R66 D<8> XDAC2/XC0/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R67 D<8> XDAC2/XC0/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R68 D<8> XDAC2/XC0/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R69 D<8> XDAC2/XC0/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R70 D<8> XDAC2/XC0/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R71 D<8> XDAC2/XC0/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R72 XA0/CN0 XDAC2/XC1/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R73 XA0/CN0 XDAC2/XC1/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R74 XA0/CN0 XDAC2/XC1/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R75 XA0/CN0 XDAC2/XC1/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R76 XA0/CN0 XDAC2/XC1/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R77 XA0/CN0 XDAC2/XC1/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R78 XA1/CN1 XDAC2/XC64b<1>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R79 XA1/CN1 XDAC2/XC64b<1>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R80 XA1/CN1 XDAC2/XC64b<1>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R81 XA1/CN1 XDAC2/XC64b<1>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R82 XA1/CN1 XDAC2/XC64b<1>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R83 XA1/CN1 XDAC2/XC64b<1>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R84 D<8> XDAC2/XC128a<1>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R85 D<8> XDAC2/XC128a<1>/XRES1A/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R86 D<8> XDAC2/XC128a<1>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R87 D<8> XDAC2/XC128a<1>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R88 D<8> XDAC2/XC128a<1>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R89 D<8> XDAC2/XC128a<1>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R90 XA2/CN1 XDAC2/XC32a<0>/XRES16/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R91 XDAC2/XC32a<0>/C1A AVSS sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R92 XA6/CN0 XDAC2/XC32a<0>/XRES2/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R93 XA7/CN0 XDAC2/XC32a<0>/XRES1B/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R94 XA5/CN0 XDAC2/XC32a<0>/XRES4/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
R95 XA4/CN0 XDAC2/XC32a<0>/XRES8/B sky130_fd_pr__res_generic_l1 w=380000u l=300000u
X0 XA20/XA9/A XA20/XA11/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.49591e+14p ps=8.019e+08u w=1.08e+06u l=180000u
X1 AVDD XA20/XA12/Y XA20/XA9/A AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X2 XA20/XA10/MN1/S XA20/XA11/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.27156e+14p ps=1.2177e+09u w=1.08e+06u l=180000u
X3 XA20/XA9/A XA20/XA12/Y XA20/XA10/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X4 XA20/XA11/MP1/S CK_SAMPLE AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X5 XA20/XA11/Y DONE XA20/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X6 XA20/XA11/Y CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X7 AVSS DONE XA20/XA11/Y AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X8 XA20/XA12/Y XA8/CEO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X9 XA20/XA12/Y XA8/CEO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X10 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X11 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X12 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X13 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X14 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X15 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X16 AVDD XA20/XA9/A XA20/XA1/MP0/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X17 XA20/XA1/MP0/S XA20/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X18 XA20/XA1/MP0/S SARP XA20/XA1/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X19 XA20/XA1/MP0/S SARP XA20/XA1/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X20 XA20/XA1/MP0/S SARP XA20/XA1/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X21 XA20/XA1/MP0/S SARP XA20/XA1/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X22 AVDD XA20/XA9/Y XA20/XA1/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=6.59084e+14p pd=1.24492e+09u as=0p ps=0u w=1.08e+06u l=180000u
X23 XA20/XA1/MP0/S SARP XA20/XA1/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X24 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X25 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X26 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X27 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X28 AVDD XA20/XA9/Y XA20/XA3/N1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X29 XA20/XA2/N2 XA20/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X30 AVDD AVDD XA20/XA2/N2 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X31 XA20/XA3/N1 XA20/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X32 XA20/XA3a/A XA20/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X33 XA20/XA2/N2 SARP XA20/XA3/N1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X34 AVDD XA20/XA3/CO XA20/XA3a/A AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X35 XA20/XA3/N1 SARP XA20/XA2/N2 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X36 XA20/XA3a/A XA20/XA3/CO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X37 XA20/XA2/N2 SARP XA20/XA3/N1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X38 AVDD XA20/XA3/CO XA20/XA3a/A AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X39 XA20/XA3/N1 SARP XA20/XA2/N2 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X40 XA20/XA3a/A XA20/XA3/CO XA20/XA2/N2 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X41 XA20/XA2/N2 SARP XA20/XA3/N1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X42 AVDD XA20/XA9/Y XA20/XA3/N1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X43 XA20/XA3/N2 XA20/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X44 AVDD AVDD XA20/XA3/N2 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X45 XA20/XA3/N1 XA20/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X46 XA20/XA3/CO XA20/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X47 XA20/XA3/N2 SARN XA20/XA3/N1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X48 AVDD XA20/XA3a/A XA20/XA3/CO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X49 XA20/XA3/N1 SARN XA20/XA3/N2 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X50 XA20/XA3/CO XA20/XA3a/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X51 XA20/XA3/N2 SARN XA20/XA3/N1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X52 AVDD XA20/XA3a/A XA20/XA3/CO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X53 XA20/XA3/N1 SARN XA20/XA3/N2 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X54 XA20/XA3/CO XA20/XA3a/A XA20/XA3/N2 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X55 XA20/XA3/N2 SARN XA20/XA3/N1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X56 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X57 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X58 AVDD XA20/XA9/A XA20/XA4/MP0/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X59 XA20/XA4/MP0/S XA20/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X60 XA20/XA4/MP0/S SARN XA20/XA4/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X61 XA20/XA4/MP0/S SARN XA20/XA4/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X62 XA20/XA4/MP0/S SARN XA20/XA4/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X63 XA20/XA4/MP0/S SARN XA20/XA4/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X64 AVDD XA20/XA9/Y XA20/XA4/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X65 XA20/XA4/MP0/S SARN XA20/XA4/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X66 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X67 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X68 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X69 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X70 XA20/CNO XA20/XA3a/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X71 AVDD XA20/XA3a/A XA20/CNO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X72 XA20/CNO XA20/XA3a/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X73 XA20/CNO XA20/XA3a/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X74 AVDD XA20/XA3a/A XA20/CNO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X75 AVSS XA20/XA3a/A XA20/CNO AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X76 XA20/CNO XA20/XA3a/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X77 AVSS XA20/XA3a/A XA20/CNO AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X78 XA20/CPO XA20/XA3/CO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X79 AVDD XA20/XA3/CO XA20/CPO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X80 XA20/CPO XA20/XA3/CO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X81 XA20/CPO XA20/XA3/CO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X82 AVDD XA20/XA3/CO XA20/CPO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X83 AVSS XA20/XA3/CO XA20/CPO AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X84 XA20/CPO XA20/XA3/CO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X85 AVSS XA20/XA3/CO XA20/CPO AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X86 XA20/XA9/Y XA20/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X87 XA20/XA9/Y XA20/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X88 SARP XB1/M4/G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=4.9248e+12p pd=2.64e+07u as=5.5404e+12p ps=2.97e+07u w=1.08e+06u l=180000u
X89 SARP XB1/M4/G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X90 SARP XB1/M4/G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X91 SARP XB1/M4/G SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X92 SARN XA0/CEIN SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=4.9248e+12p pd=2.64e+07u as=0p ps=0u w=1.08e+06u l=180000u
R96 XB1/XA4/GNG XB1/XCAPB1/XCAPB0/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R97 XB1/XCAPB1/XCAPB0/m3_252_308# XB1/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R98 XB1/XA4/GNG XB1/XCAPB1/XCAPB1/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R99 XB1/XCAPB1/XCAPB1/m3_252_308# XB1/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R100 XB1/XA4/GNG XB1/XCAPB1/XCAPB2/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R101 XB1/XCAPB1/XCAPB2/m3_252_308# XB1/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R102 XB1/XA4/GNG XB1/XCAPB1/XCAPB3/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R103 XB1/XCAPB1/XCAPB3/m3_252_308# XB1/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R104 XB1/XA4/GNG XB1/XCAPB1/XCAPB4/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R105 XB1/XCAPB1/XCAPB4/m3_252_308# XB1/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
X93 SARN XA0/CEIN SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X94 SARN XA0/CEIN SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X95 SARN XA0/CEIN SAR_IP AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X96 XB1/CKN CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X97 XB1/CKN CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X98 XB1/XA1/Y XB1/XA1/MP0/G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X99 XB1/XA1/MP0/G XB1/XA1/MP0/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X100 XB1/XA2/MP0/G XB1/XA2/MP0/G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X101 XA0/CEIN XB1/XA2/MP0/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X102 XB1/XA3/B AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X103 AVDD XB1/CKN XB1/XA3/MP0/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X104 SAR_IP XB1/CKN XB1/XA3/B AVDD sky130_fd_pr__pfet_01v8 ad=6.156e+11p pd=3.3e+06u as=0p ps=0u w=1.08e+06u l=180000u
X105 AVSS XB1/CKN XB1/XA3/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X106 XB1/XA3/B XB1/CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X107 SAR_IP XB1/XA3/MP0/S XB1/XA3/B AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X108 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X109 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X110 XB1/XA4/GNG XB1/CKN XB1/M4/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X111 AVDD XB1/M4/G XB1/XA4/GNG AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X112 XB1/XA4/MN1/S XB1/CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X113 XB1/M4/G XB1/XA1/Y XB1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X114 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X115 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X116 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X117 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X118 XA0/XA11/A XA0/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X119 XA0/XA11/A XA0/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X120 XA0/XA11/MP1/S XA0/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X121 XA0/XA12/A XA0/CEIN XA0/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X122 XA0/XA12/A XA0/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X123 AVSS XA0/CEIN XA0/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X124 XA0/CEO XA0/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X125 XA0/CEO XA0/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X126 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X127 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X128 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X129 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X130 AVDD EN XA0/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X131 XA0/XA1/XA1/MP2/S XA20/CNO XA1/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X132 XA0/XA1/XA1/MP3/S XA20/CPO XA0/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X133 XA0/XA1/XA1/MN2/S EN XA0/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X134 AVDD XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X135 XA0/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X136 AVSS XA20/CPO XA0/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X137 XA1/EN XA0/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X138 XA0/XA1/XA2/Y XA1/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X139 XA0/XA1/XA2/Y XA1/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X140 XA0/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X141 XA0/XA1/XA4/MP2/S EN XA0/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X142 XA0/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X143 XA0/XA4/A EN XA0/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X144 XA0/XA1/XA4/MN2/S XA0/XA1/XA2/Y XA0/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X145 XA0/XA4/A EN XA0/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X146 XA0/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X147 XA0/XA1/XA5/MP2/S EN XA0/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X148 XA0/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X149 XA0/XA2/A EN XA0/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X150 XA0/XA1/XA5/MN2/S XA0/XA1/XA2/Y XA0/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X151 XA0/XA2/A EN XA0/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X152 D<8> XA0/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=8.86464e+13p ps=4.752e+08u w=1.08e+06u l=180000u
X153 VREF XA0/XA2/A D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X154 D<8> XA0/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X155 D<8> XA0/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X156 VREF XA0/XA2/A D<8> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X157 AVSS XA0/XA2/A D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X158 D<8> XA0/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X159 AVSS XA0/XA2/A D<8> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X160 XA0/CP1 D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X161 VREF D<8> XA0/CP1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X162 XA0/CP1 D<8> VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X163 XA0/CP1 D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X164 VREF D<8> XA0/CP1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X165 AVSS D<8> XA0/CP1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X166 XA0/CP1 D<8> AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X167 AVSS D<8> XA0/CP1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X168 XA0/CP0 XA0/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X169 VREF XA0/XA4/A XA0/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X170 XA0/CP0 XA0/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X171 XA0/CP0 XA0/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X172 VREF XA0/XA4/A XA0/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X173 AVSS XA0/XA4/A XA0/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X174 XA0/CP0 XA0/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X175 AVSS XA0/XA4/A XA0/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X176 XA0/CN0 XA0/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X177 VREF XA0/CP0 XA0/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X178 XA0/CN0 XA0/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X179 XA0/CN0 XA0/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X180 VREF XA0/CP0 XA0/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X181 AVSS XA0/CP0 XA0/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X182 XA0/CN0 XA0/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X183 AVSS XA0/CP0 XA0/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X184 XA0/XA6/MP1/S XA0/CN0 XA0/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X185 AVDD XA0/CN0 XA0/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X186 XA0/XA6/MP3/S XA0/CP1 AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X187 XA0/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X188 XA0/XA9/B XA0/CP1 XA0/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X189 AVSS CK_SAMPLE XA0/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X190 XA0/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X191 XA0/XA9/B CK_SAMPLE XA0/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X192 XA0/XA9/A XA1/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X193 XA0/XA9/A XA1/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X194 XA0/DONE XA0/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X195 XA0/DONE XA0/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X196 XA0/XA9/Y XA0/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X197 AVDD XA0/XA9/B XA0/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X198 XA0/XA9/MN1/S XA0/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X199 XA0/XA9/Y XA0/XA9/B XA0/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X200 SARN XB2/M4/G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.5404e+12p ps=2.97e+07u w=1.08e+06u l=180000u
X201 SARN XB2/M4/G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X202 SARN XB2/M4/G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X203 SARN XB2/M4/G SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X204 SARP XA0/CEIN SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
R106 XB2/XA4/GNG XB2/XCAPB1/XCAPB0/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R107 XB2/XCAPB1/XCAPB0/m3_252_308# XB2/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R108 XB2/XA4/GNG XB2/XCAPB1/XCAPB1/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R109 XB2/XCAPB1/XCAPB1/m3_252_308# XB2/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R110 XB2/XA4/GNG XB2/XCAPB1/XCAPB2/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R111 XB2/XCAPB1/XCAPB2/m3_252_308# XB2/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R112 XB2/XA4/GNG XB2/XCAPB1/XCAPB3/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R113 XB2/XCAPB1/XCAPB3/m3_252_308# XB2/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R114 XB2/XA4/GNG XB2/XCAPB1/XCAPB4/m3_9828_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R115 XB2/XCAPB1/XCAPB4/m3_252_308# XB2/XA3/B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
X205 SARP XA0/CEIN SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X206 SARP XA0/CEIN SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X207 SARP XA0/CEIN SAR_IN AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X208 XB2/CKN CK_SAMPLE_BSSW AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X209 XB2/CKN CK_SAMPLE_BSSW AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X210 XB2/XA1/Y XB2/XA1/MP0/G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X211 XB2/XA1/MP0/G XB2/XA1/MP0/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X212 XB2/XA2/MP0/G XB2/XA2/MP0/G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X213 XA0/CEIN XB2/XA2/MP0/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X214 XB2/XA3/B AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X215 AVDD XB2/CKN XB2/XA3/MP0/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X216 SAR_IN XB2/CKN XB2/XA3/B AVDD sky130_fd_pr__pfet_01v8 ad=6.156e+11p pd=3.3e+06u as=0p ps=0u w=1.08e+06u l=180000u
X217 AVSS XB2/CKN XB2/XA3/MP0/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X218 XB2/XA3/B XB2/CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X219 SAR_IN XB2/XA3/MP0/S XB2/XA3/B AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X220 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X221 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X222 XB2/XA4/GNG XB2/CKN XB2/M4/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X223 AVDD XB2/M4/G XB2/XA4/GNG AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X224 XB2/XA4/MN1/S XB2/CKN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X225 XB2/M4/G XB2/XA1/Y XB2/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X226 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X227 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X228 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X229 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X230 XA1/XA11/A XA1/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X231 XA1/XA11/A XA1/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X232 XA1/XA11/MP1/S XA1/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X233 XA1/XA12/A XA0/CEO XA1/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X234 XA1/XA12/A XA1/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X235 AVSS XA0/CEO XA1/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X236 XA1/CEO XA1/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X237 XA1/CEO XA1/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X239 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X240 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X241 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X242 AVDD EN XA1/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X243 XA1/XA1/XA1/MP2/S XA20/CNO XA2/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X244 XA1/XA1/XA1/MP3/S XA20/CPO XA1/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X245 XA1/XA1/XA1/MN2/S XA1/EN XA1/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X246 AVDD XA1/XA1/XA1/MP3/G XA1/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X247 XA1/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X248 AVSS XA20/CPO XA1/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X249 XA2/EN XA1/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X250 XA1/XA1/XA2/Y XA2/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X251 XA1/XA1/XA2/Y XA2/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X252 XA1/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X253 XA1/XA1/XA4/MP2/S EN XA1/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X254 XA1/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X255 XA1/XA4/A EN XA1/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X256 XA1/XA1/XA4/MN2/S XA1/XA1/XA2/Y XA1/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X257 XA1/XA4/A XA1/EN XA1/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X258 XA1/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X259 XA1/XA1/XA5/MP2/S EN XA1/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X260 XA1/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X261 XA1/XA2/A EN XA1/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X262 XA1/XA1/XA5/MN2/S XA1/XA1/XA2/Y XA1/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X263 XA1/XA2/A XA1/EN XA1/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X264 XA1/CN1 XA1/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X265 VREF XA1/XA2/A XA1/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X266 XA1/CN1 XA1/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X267 XA1/CN1 XA1/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X268 VREF XA1/XA2/A XA1/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X269 AVSS XA1/XA2/A XA1/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X270 XA1/CN1 XA1/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X271 AVSS XA1/XA2/A XA1/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X272 D<7> XA1/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X273 VREF XA1/CN1 D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X274 D<7> XA1/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X275 D<7> XA1/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X276 VREF XA1/CN1 D<7> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X277 AVSS XA1/CN1 D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X278 D<7> XA1/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X279 AVSS XA1/CN1 D<7> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X280 XA1/CP0 XA1/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X281 VREF XA1/XA4/A XA1/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X282 XA1/CP0 XA1/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X283 XA1/CP0 XA1/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X284 VREF XA1/XA4/A XA1/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X285 AVSS XA1/XA4/A XA1/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X286 XA1/CP0 XA1/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X287 AVSS XA1/XA4/A XA1/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X288 XA1/CN0 XA1/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X289 VREF XA1/CP0 XA1/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X290 XA1/CN0 XA1/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X291 XA1/CN0 XA1/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X292 VREF XA1/CP0 XA1/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X293 AVSS XA1/CP0 XA1/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X294 XA1/CN0 XA1/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X295 AVSS XA1/CP0 XA1/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X296 XA1/XA6/MP1/S XA1/CN0 XA1/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X297 AVDD XA1/CN0 XA1/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X298 XA1/XA6/MP3/S D<7> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X299 XA1/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X300 XA1/XA9/B D<7> XA1/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X301 AVSS CK_SAMPLE XA1/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X302 XA1/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X303 XA1/XA9/B CK_SAMPLE XA1/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X304 XA1/XA9/A XA2/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X305 XA1/XA9/A XA2/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X306 XA1/DONE XA1/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X307 XA1/DONE XA1/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X308 XA1/XA9/Y XA1/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X309 AVDD XA1/XA9/B XA1/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X310 XA1/XA9/MN1/S XA1/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X311 XA1/XA9/Y XA1/XA9/B XA1/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X312 XA2/XA11/A XA2/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X313 XA2/XA11/A XA2/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X314 XA2/XA11/MP1/S XA2/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X315 XA2/XA12/A XA1/CEO XA2/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X316 XA2/XA12/A XA2/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X317 AVSS XA1/CEO XA2/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X318 XA2/CEO XA2/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X319 XA2/CEO XA2/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X320 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X321 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X322 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X323 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X324 AVDD EN XA2/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X325 XA2/XA1/XA1/MP2/S XA20/CNO XA3/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X326 XA2/XA1/XA1/MP3/S XA20/CPO XA2/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X327 XA2/XA1/XA1/MN2/S XA2/EN XA2/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X328 AVDD XA2/XA1/XA1/MP3/G XA2/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X329 XA2/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X330 AVSS XA20/CPO XA2/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X331 XA3/EN XA2/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X332 XA2/XA1/XA2/Y XA3/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X333 XA2/XA1/XA2/Y XA3/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X334 XA2/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X335 XA2/XA1/XA4/MP2/S EN XA2/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X336 XA2/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X337 XA2/XA4/A EN XA2/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X338 XA2/XA1/XA4/MN2/S XA2/XA1/XA2/Y XA2/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X339 XA2/XA4/A XA2/EN XA2/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X340 XA2/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X341 XA2/XA1/XA5/MP2/S EN XA2/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X342 XA2/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X343 XA2/XA2/A EN XA2/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X344 XA2/XA1/XA5/MN2/S XA2/XA1/XA2/Y XA2/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X345 XA2/XA2/A XA2/EN XA2/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X346 XA2/CN1 XA2/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X347 VREF XA2/XA2/A XA2/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X348 XA2/CN1 XA2/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X349 XA2/CN1 XA2/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X350 VREF XA2/XA2/A XA2/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X351 AVSS XA2/XA2/A XA2/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X352 XA2/CN1 XA2/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X353 AVSS XA2/XA2/A XA2/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X354 D<6> XA2/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X355 VREF XA2/CN1 D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X356 D<6> XA2/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X357 D<6> XA2/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X358 VREF XA2/CN1 D<6> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X359 AVSS XA2/CN1 D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X360 D<6> XA2/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X361 AVSS XA2/CN1 D<6> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X362 XA2/CP0 XA2/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X363 VREF XA2/XA4/A XA2/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X364 XA2/CP0 XA2/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X365 XA2/CP0 XA2/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X366 VREF XA2/XA4/A XA2/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X367 AVSS XA2/XA4/A XA2/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X368 XA2/CP0 XA2/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X369 AVSS XA2/XA4/A XA2/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X370 XA2/CN0 XA2/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X371 VREF XA2/CP0 XA2/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X372 XA2/CN0 XA2/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X373 XA2/CN0 XA2/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X374 VREF XA2/CP0 XA2/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X375 AVSS XA2/CP0 XA2/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X376 XA2/CN0 XA2/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X377 AVSS XA2/CP0 XA2/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X378 XA2/XA6/MP1/S XA2/CN0 XA2/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X379 AVDD XA2/CN0 XA2/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X380 XA2/XA6/MP3/S D<6> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X381 XA2/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X382 XA2/XA9/B D<6> XA2/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X383 AVSS CK_SAMPLE XA2/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X384 XA2/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X385 XA2/XA9/B CK_SAMPLE XA2/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X386 XA2/XA9/A XA3/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X387 XA2/XA9/A XA3/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X388 XA2/DONE XA2/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X389 XA2/DONE XA2/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X390 XA2/XA9/Y XA2/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X391 AVDD XA2/XA9/B XA2/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X392 XA2/XA9/MN1/S XA2/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X393 XA2/XA9/Y XA2/XA9/B XA2/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X394 XA3/XA11/A XA3/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X395 XA3/XA11/A XA3/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X396 XA3/XA11/MP1/S XA3/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X397 XA3/XA12/A XA2/CEO XA3/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X398 XA3/XA12/A XA3/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X399 AVSS XA2/CEO XA3/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X400 XA3/CEO XA3/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X401 XA3/CEO XA3/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X402 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X403 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X404 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X405 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X406 AVDD EN XA3/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X407 XA3/XA1/XA1/MP2/S XA20/CNO XA4/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X408 XA3/XA1/XA1/MP3/S XA20/CPO XA3/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X409 XA3/XA1/XA1/MN2/S XA3/EN XA3/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X410 AVDD XA3/XA1/XA1/MP3/G XA3/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X411 XA3/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X412 AVSS XA20/CPO XA3/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X413 XA4/EN XA3/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X414 XA3/XA1/XA2/Y XA4/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X415 XA3/XA1/XA2/Y XA4/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X416 XA3/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X417 XA3/XA1/XA4/MP2/S EN XA3/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X418 XA3/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X419 XA3/XA4/A EN XA3/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X420 XA3/XA1/XA4/MN2/S XA3/XA1/XA2/Y XA3/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X421 XA3/XA4/A XA3/EN XA3/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X422 XA3/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X423 XA3/XA1/XA5/MP2/S EN XA3/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X424 XA3/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X425 XA3/XA2/A EN XA3/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X426 XA3/XA1/XA5/MN2/S XA3/XA1/XA2/Y XA3/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X427 XA3/XA2/A XA3/EN XA3/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X428 XA3/CN1 XA3/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X429 VREF XA3/XA2/A XA3/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X430 XA3/CN1 XA3/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X431 XA3/CN1 XA3/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X432 VREF XA3/XA2/A XA3/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X433 AVSS XA3/XA2/A XA3/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X434 XA3/CN1 XA3/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X435 AVSS XA3/XA2/A XA3/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X436 D<5> XA3/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X437 VREF XA3/CN1 D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X438 D<5> XA3/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X439 D<5> XA3/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X440 VREF XA3/CN1 D<5> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X441 AVSS XA3/CN1 D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X442 D<5> XA3/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X443 AVSS XA3/CN1 D<5> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X444 XA3/CP0 XA3/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X445 VREF XA3/XA4/A XA3/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X446 XA3/CP0 XA3/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X447 XA3/CP0 XA3/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X448 VREF XA3/XA4/A XA3/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X449 AVSS XA3/XA4/A XA3/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X450 XA3/CP0 XA3/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X451 AVSS XA3/XA4/A XA3/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X452 XA3/CN0 XA3/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X453 VREF XA3/CP0 XA3/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X454 XA3/CN0 XA3/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X455 XA3/CN0 XA3/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X456 VREF XA3/CP0 XA3/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X457 AVSS XA3/CP0 XA3/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X458 XA3/CN0 XA3/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X459 AVSS XA3/CP0 XA3/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X460 XA3/XA6/MP1/S XA3/CN0 XA3/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X461 AVDD XA3/CN0 XA3/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X462 XA3/XA6/MP3/S D<5> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X463 XA3/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X464 XA3/XA9/B D<5> XA3/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X465 AVSS CK_SAMPLE XA3/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X466 XA3/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X467 XA3/XA9/B CK_SAMPLE XA3/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X468 XA3/XA9/A XA4/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X469 XA3/XA9/A XA4/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X470 XA3/DONE XA3/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X471 XA3/DONE XA3/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X472 XA3/XA9/Y XA3/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X473 AVDD XA3/XA9/B XA3/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X474 XA3/XA9/MN1/S XA3/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X475 XA3/XA9/Y XA3/XA9/B XA3/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X476 XA4/XA11/A XA4/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X477 XA4/XA11/A XA4/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X478 XA4/XA11/MP1/S XA4/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X479 XA4/XA12/A XA3/CEO XA4/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X480 XA4/XA12/A XA4/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X481 AVSS XA3/CEO XA4/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X482 XA4/CEO XA4/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X483 XA4/CEO XA4/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X484 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X485 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X486 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X487 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X488 AVDD EN XA4/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X489 XA4/XA1/XA1/MP2/S XA20/CNO XA5/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X490 XA4/XA1/XA1/MP3/S XA20/CPO XA4/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X491 XA4/XA1/XA1/MN2/S XA4/EN XA4/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X492 AVDD XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X493 XA4/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X494 AVSS XA20/CPO XA4/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X495 XA5/EN XA4/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X496 XA4/XA1/XA2/Y XA5/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X497 XA4/XA1/XA2/Y XA5/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X498 XA4/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X499 XA4/XA1/XA4/MP2/S EN XA4/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X500 XA4/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X501 XA4/XA4/A EN XA4/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X502 XA4/XA1/XA4/MN2/S XA4/XA1/XA2/Y XA4/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X503 XA4/XA4/A XA4/EN XA4/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X504 XA4/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X505 XA4/XA1/XA5/MP2/S EN XA4/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X506 XA4/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X507 XA4/XA2/A EN XA4/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X508 XA4/XA1/XA5/MN2/S XA4/XA1/XA2/Y XA4/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X509 XA4/XA2/A XA4/EN XA4/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X510 XA4/CN1 XA4/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X511 VREF XA4/XA2/A XA4/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X512 XA4/CN1 XA4/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X513 XA4/CN1 XA4/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X514 VREF XA4/XA2/A XA4/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X515 AVSS XA4/XA2/A XA4/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X516 XA4/CN1 XA4/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X517 AVSS XA4/XA2/A XA4/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X518 D<4> XA4/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X519 VREF XA4/CN1 D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X520 D<4> XA4/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X521 D<4> XA4/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X522 VREF XA4/CN1 D<4> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X523 AVSS XA4/CN1 D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X524 D<4> XA4/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X525 AVSS XA4/CN1 D<4> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X526 XA4/CP0 XA4/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X527 VREF XA4/XA4/A XA4/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X528 XA4/CP0 XA4/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X529 XA4/CP0 XA4/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X530 VREF XA4/XA4/A XA4/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X531 AVSS XA4/XA4/A XA4/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X532 XA4/CP0 XA4/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X533 AVSS XA4/XA4/A XA4/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X534 XA4/CN0 XA4/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X535 VREF XA4/CP0 XA4/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X536 XA4/CN0 XA4/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X537 XA4/CN0 XA4/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X538 VREF XA4/CP0 XA4/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X539 AVSS XA4/CP0 XA4/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X540 XA4/CN0 XA4/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X541 AVSS XA4/CP0 XA4/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X542 XA4/XA6/MP1/S XA4/CN0 XA4/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X543 AVDD XA4/CN0 XA4/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X544 XA4/XA6/MP3/S D<4> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X545 XA4/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X546 XA4/XA9/B D<4> XA4/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X547 AVSS CK_SAMPLE XA4/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X548 XA4/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X549 XA4/XA9/B CK_SAMPLE XA4/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X550 XA4/XA9/A XA5/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X551 XA4/XA9/A XA5/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X552 XA4/DONE XA4/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X553 XA4/DONE XA4/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X554 XA4/XA9/Y XA4/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X555 AVDD XA4/XA9/B XA4/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X556 XA4/XA9/MN1/S XA4/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X557 XA4/XA9/Y XA4/XA9/B XA4/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X558 XA5/XA11/A XA5/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X559 XA5/XA11/A XA5/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X560 XA5/XA11/MP1/S XA5/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X561 XA5/XA12/A XA4/CEO XA5/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X562 XA5/XA12/A XA5/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X563 AVSS XA4/CEO XA5/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X564 XA5/CEO XA5/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X565 XA5/CEO XA5/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X566 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X567 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X568 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X569 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X570 AVDD EN XA5/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X571 XA5/XA1/XA1/MP2/S XA20/CNO XA6/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X572 XA5/XA1/XA1/MP3/S XA20/CPO XA5/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X573 XA5/XA1/XA1/MN2/S XA5/EN XA5/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X574 AVDD XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X575 XA5/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X576 AVSS XA20/CPO XA5/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X577 XA6/EN XA5/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X578 XA5/XA1/XA2/Y XA6/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X579 XA5/XA1/XA2/Y XA6/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X580 XA5/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X581 XA5/XA1/XA4/MP2/S EN XA5/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X582 XA5/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X583 XA5/XA4/A EN XA5/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X584 XA5/XA1/XA4/MN2/S XA5/XA1/XA2/Y XA5/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X585 XA5/XA4/A XA5/EN XA5/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X586 XA5/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X587 XA5/XA1/XA5/MP2/S EN XA5/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X588 XA5/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X589 XA5/XA2/A EN XA5/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X590 XA5/XA1/XA5/MN2/S XA5/XA1/XA2/Y XA5/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X591 XA5/XA2/A XA5/EN XA5/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X592 XA5/CN1 XA5/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X593 VREF XA5/XA2/A XA5/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X594 XA5/CN1 XA5/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X595 XA5/CN1 XA5/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X596 VREF XA5/XA2/A XA5/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X597 AVSS XA5/XA2/A XA5/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X598 XA5/CN1 XA5/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X599 AVSS XA5/XA2/A XA5/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X600 D<3> XA5/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X601 VREF XA5/CN1 D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X602 D<3> XA5/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X603 D<3> XA5/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X604 VREF XA5/CN1 D<3> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X605 AVSS XA5/CN1 D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X606 D<3> XA5/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X607 AVSS XA5/CN1 D<3> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X608 XA5/CP0 XA5/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X609 VREF XA5/XA4/A XA5/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X610 XA5/CP0 XA5/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X611 XA5/CP0 XA5/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X612 VREF XA5/XA4/A XA5/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X613 AVSS XA5/XA4/A XA5/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X614 XA5/CP0 XA5/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X615 AVSS XA5/XA4/A XA5/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X616 XA5/CN0 XA5/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X617 VREF XA5/CP0 XA5/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X618 XA5/CN0 XA5/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X619 XA5/CN0 XA5/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X620 VREF XA5/CP0 XA5/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X621 AVSS XA5/CP0 XA5/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X622 XA5/CN0 XA5/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X623 AVSS XA5/CP0 XA5/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X624 XA5/XA6/MP1/S XA5/CN0 XA5/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X625 AVDD XA5/CN0 XA5/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X626 XA5/XA6/MP3/S D<3> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X627 XA5/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X628 XA5/XA9/B D<3> XA5/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X629 AVSS CK_SAMPLE XA5/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X630 XA5/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X631 XA5/XA9/B CK_SAMPLE XA5/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X632 XA5/XA9/A XA6/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X633 XA5/XA9/A XA6/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X634 XA5/DONE XA5/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X635 XA5/DONE XA5/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X636 XA5/XA9/Y XA5/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X637 AVDD XA5/XA9/B XA5/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X638 XA5/XA9/MN1/S XA5/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X639 XA5/XA9/Y XA5/XA9/B XA5/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X640 XA6/XA11/A XA6/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X641 XA6/XA11/A XA6/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X642 XA6/XA11/MP1/S XA6/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X643 XA6/XA12/A XA5/CEO XA6/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X644 XA6/XA12/A XA6/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X645 AVSS XA5/CEO XA6/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X646 XA6/CEO XA6/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X647 XA6/CEO XA6/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X648 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X649 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X650 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X651 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X652 AVDD EN XA6/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X653 XA6/XA1/XA1/MP2/S XA20/CNO XA7/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X654 XA6/XA1/XA1/MP3/S XA20/CPO XA6/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X655 XA6/XA1/XA1/MN2/S XA6/EN XA6/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X656 AVDD XA6/XA1/XA1/MP3/G XA6/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X657 XA6/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X658 AVSS XA20/CPO XA6/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X659 XA7/EN XA6/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X660 XA6/XA1/XA2/Y XA7/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X661 XA6/XA1/XA2/Y XA7/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X662 XA6/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X663 XA6/XA1/XA4/MP2/S EN XA6/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X664 XA6/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X665 XA6/XA4/A EN XA6/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X666 XA6/XA1/XA4/MN2/S XA6/XA1/XA2/Y XA6/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X667 XA6/XA4/A XA6/EN XA6/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X668 XA6/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X669 XA6/XA1/XA5/MP2/S EN XA6/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X670 XA6/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X671 XA6/XA2/A EN XA6/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X672 XA6/XA1/XA5/MN2/S XA6/XA1/XA2/Y XA6/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X673 XA6/XA2/A XA6/EN XA6/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X674 XA6/CN1 XA6/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X675 VREF XA6/XA2/A XA6/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X676 XA6/CN1 XA6/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X677 XA6/CN1 XA6/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X678 VREF XA6/XA2/A XA6/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X679 AVSS XA6/XA2/A XA6/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X680 XA6/CN1 XA6/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X681 AVSS XA6/XA2/A XA6/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X682 D<2> XA6/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X683 VREF XA6/CN1 D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X684 D<2> XA6/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X685 D<2> XA6/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X686 VREF XA6/CN1 D<2> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X687 AVSS XA6/CN1 D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X688 D<2> XA6/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X689 AVSS XA6/CN1 D<2> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X690 XA6/CP0 XA6/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X691 VREF XA6/XA4/A XA6/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X692 XA6/CP0 XA6/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X693 XA6/CP0 XA6/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X694 VREF XA6/XA4/A XA6/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X695 AVSS XA6/XA4/A XA6/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X696 XA6/CP0 XA6/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X697 AVSS XA6/XA4/A XA6/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X698 XA6/CN0 XA6/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X699 VREF XA6/CP0 XA6/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X700 XA6/CN0 XA6/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X701 XA6/CN0 XA6/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X702 VREF XA6/CP0 XA6/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X703 AVSS XA6/CP0 XA6/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X704 XA6/CN0 XA6/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X705 AVSS XA6/CP0 XA6/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X706 XA6/XA6/MP1/S XA6/CN0 XA6/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X707 AVDD XA6/CN0 XA6/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X708 XA6/XA6/MP3/S D<2> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X709 XA6/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X710 XA6/XA9/B D<2> XA6/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X711 AVSS CK_SAMPLE XA6/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X712 XA6/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X713 XA6/XA9/B CK_SAMPLE XA6/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X714 XA6/XA9/A XA7/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X715 XA6/XA9/A XA7/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X716 XA6/DONE XA6/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X717 XA6/DONE XA6/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X718 XA6/XA9/Y XA6/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X719 AVDD XA6/XA9/B XA6/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X720 XA6/XA9/MN1/S XA6/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X721 XA6/XA9/Y XA6/XA9/B XA6/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X722 XA7/XA11/A XA7/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X723 XA7/XA11/A XA7/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X724 XA7/XA11/MP1/S XA7/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X725 XA7/XA12/A XA6/CEO XA7/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X726 XA7/XA12/A XA7/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X727 AVSS XA6/CEO XA7/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X728 XA7/CEO XA7/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X729 XA7/CEO XA7/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X730 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X731 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X732 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X733 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X734 AVDD EN XA7/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X735 XA7/XA1/XA1/MP2/S XA20/CNO XA8/EN AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X736 XA7/XA1/XA1/MP3/S XA20/CPO XA7/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X737 XA7/XA1/XA1/MN2/S XA7/EN XA7/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X738 AVDD XA7/XA1/XA1/MP3/G XA7/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X739 XA7/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X740 AVSS XA20/CPO XA7/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X741 XA8/EN XA7/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X742 XA7/XA1/XA2/Y XA8/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X743 XA7/XA1/XA2/Y XA8/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X744 XA7/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X745 XA7/XA1/XA4/MP2/S EN XA7/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X746 XA7/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X747 XA7/XA4/A EN XA7/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X748 XA7/XA1/XA4/MN2/S XA7/XA1/XA2/Y XA7/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X749 XA7/XA4/A XA7/EN XA7/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X750 XA7/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X751 XA7/XA1/XA5/MP2/S EN XA7/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X752 XA7/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X753 XA7/XA2/A EN XA7/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X754 XA7/XA1/XA5/MN2/S XA7/XA1/XA2/Y XA7/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X755 XA7/XA2/A XA7/EN XA7/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X756 XA7/CN1 XA7/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X757 VREF XA7/XA2/A XA7/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X758 XA7/CN1 XA7/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X759 XA7/CN1 XA7/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X760 VREF XA7/XA2/A XA7/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X761 AVSS XA7/XA2/A XA7/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X762 XA7/CN1 XA7/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X763 AVSS XA7/XA2/A XA7/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X764 D<1> XA7/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X765 VREF XA7/CN1 D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X766 D<1> XA7/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X767 D<1> XA7/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X768 VREF XA7/CN1 D<1> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X769 AVSS XA7/CN1 D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X770 D<1> XA7/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X771 AVSS XA7/CN1 D<1> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X772 XA7/CP0 XA7/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X773 VREF XA7/XA4/A XA7/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X774 XA7/CP0 XA7/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X775 XA7/CP0 XA7/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X776 VREF XA7/XA4/A XA7/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X777 AVSS XA7/XA4/A XA7/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X778 XA7/CP0 XA7/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X779 AVSS XA7/XA4/A XA7/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X780 XA7/CN0 XA7/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X781 VREF XA7/CP0 XA7/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X782 XA7/CN0 XA7/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X783 XA7/CN0 XA7/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X784 VREF XA7/CP0 XA7/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X785 AVSS XA7/CP0 XA7/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X786 XA7/CN0 XA7/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X787 AVSS XA7/CP0 XA7/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X788 XA7/XA6/MP1/S XA7/CN0 XA7/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X789 AVDD XA7/CN0 XA7/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X790 XA7/XA6/MP3/S D<1> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X791 XA7/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X792 XA7/XA9/B D<1> XA7/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X793 AVSS CK_SAMPLE XA7/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X794 XA7/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X795 XA7/XA9/B CK_SAMPLE XA7/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X796 XA7/XA9/A XA8/EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X797 XA7/XA9/A XA8/EN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X798 XA7/DONE XA7/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X799 XA7/DONE XA7/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X800 XA7/XA9/Y XA7/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X801 AVDD XA7/XA9/B XA7/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X802 XA7/XA9/MN1/S XA7/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X803 XA7/XA9/Y XA7/XA9/B XA7/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X804 XA8/XA11/A XA8/XA9/Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X805 XA8/XA11/A XA8/XA9/Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X806 XA8/XA11/MP1/S XA8/XA11/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X807 XA8/XA12/A XA7/CEO XA8/XA11/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X808 XA8/XA12/A XA8/XA11/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X809 AVSS XA7/CEO XA8/XA12/A AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X810 XA8/CEO XA8/XA12/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X811 XA8/CEO XA8/XA12/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X812 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X813 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X814 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X815 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X816 AVDD EN XA8/XA1/XA1/MP3/G AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X817 XA8/XA1/XA1/MP2/S XA20/CNO XA8/ENO AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X818 XA8/XA1/XA1/MP3/S XA20/CPO XA8/XA1/XA1/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X819 XA8/XA1/XA1/MN2/S XA8/EN XA8/XA1/XA1/MP3/G AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X820 AVDD XA8/XA1/XA1/MP3/G XA8/XA1/XA1/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X821 XA8/XA1/XA1/MN2/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X822 AVSS XA20/CPO XA8/XA1/XA1/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X823 XA8/ENO XA8/XA1/XA1/MP3/G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X824 XA8/XA1/XA2/Y XA8/ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X825 XA8/XA1/XA2/Y XA8/ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X826 XA8/XA1/XA4/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X827 XA8/XA1/XA4/MP2/S EN XA8/XA1/XA4/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X828 XA8/XA1/XA4/MN1/S XA20/CPO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X829 XA8/XA4/A EN XA8/XA1/XA4/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X830 XA8/XA1/XA4/MN2/S XA8/XA1/XA2/Y XA8/XA1/XA4/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X831 XA8/XA4/A XA8/EN XA8/XA1/XA4/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X832 XA8/XA1/XA5/MP1/S EN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X833 XA8/XA1/XA5/MP2/S EN XA8/XA1/XA5/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X834 XA8/XA1/XA5/MN1/S XA20/CNO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X835 XA8/XA2/A EN XA8/XA1/XA5/MP2/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X836 XA8/XA1/XA5/MN2/S XA8/XA1/XA2/Y XA8/XA1/XA5/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X837 XA8/XA2/A XA8/EN XA8/XA1/XA5/MN2/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X838 XA8/CN1 XA8/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X839 VREF XA8/XA2/A XA8/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X840 XA8/CN1 XA8/XA2/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X841 XA8/CN1 XA8/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X842 VREF XA8/XA2/A XA8/CN1 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X843 AVSS XA8/XA2/A XA8/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X844 XA8/CN1 XA8/XA2/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X845 AVSS XA8/XA2/A XA8/CN1 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X846 D<0> XA8/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X847 VREF XA8/CN1 D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X848 D<0> XA8/CN1 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X849 D<0> XA8/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X850 VREF XA8/CN1 D<0> AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X851 AVSS XA8/CN1 D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X852 D<0> XA8/CN1 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X853 AVSS XA8/CN1 D<0> AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X854 XA8/CP0 XA8/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X855 VREF XA8/XA4/A XA8/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X856 XA8/CP0 XA8/XA4/A VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X857 XA8/CP0 XA8/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X858 VREF XA8/XA4/A XA8/CP0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X859 AVSS XA8/XA4/A XA8/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X860 XA8/CP0 XA8/XA4/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X861 AVSS XA8/XA4/A XA8/CP0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X862 XA8/CN0 XA8/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X863 VREF XA8/CP0 XA8/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X864 XA8/CN0 XA8/CP0 VREF AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X865 XA8/CN0 XA8/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X866 VREF XA8/CP0 XA8/CN0 AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X867 AVSS XA8/CP0 XA8/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X868 XA8/CN0 XA8/CP0 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X869 AVSS XA8/CP0 XA8/CN0 AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X870 XA8/XA6/MP1/S XA8/CN0 XA8/XA9/B AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X871 AVDD XA8/CN0 XA8/XA6/MP1/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X872 XA8/XA6/MP3/S D<0> AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X873 XA8/XA6/MN1/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X874 XA8/XA9/B D<0> XA8/XA6/MP3/S AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X875 AVSS CK_SAMPLE XA8/XA6/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X876 XA8/XA6/MN3/S CK_SAMPLE AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X877 XA8/XA9/B CK_SAMPLE XA8/XA6/MN3/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X878 XA8/XA9/A XA8/ENO AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X879 XA8/XA9/A XA8/ENO AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X880 DONE XA8/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=6.156e+11p pd=3.3e+06u as=0p ps=0u w=1.08e+06u l=180000u
X881 DONE XA8/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=6.156e+11p pd=3.3e+06u as=0p ps=0u w=1.08e+06u l=180000u
X882 XA8/XA9/Y XA8/XA9/A AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X883 AVDD XA8/XA9/B XA8/XA9/Y AVDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X884 XA8/XA9/MN1/S XA8/XA9/A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X885 XA8/XA9/Y XA8/XA9/B XA8/XA9/MN1/S AVSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
C0 XDAC2/XC64a<0>/XRES16/B XA0/CN0 0.05fF
C1 D<2> XDAC1/XC32a<0>/XRES16/B 0.02fF
C2 XA7/XA5/MP0/a_216_n18# VREF 0.02fF
C3 XA7/XA5/MP1/a_216_n18# VREF 0.02fF
C4 XDAC1/XC64a<0>/XRES4/B XDAC1/XC64a<0>/XRES2/B 0.55fF
C5 XA2/XA8/MP0/a_216_n18# XA3/EN 0.08fF
C6 XDAC1/XC128a<1>/XRES16/B AVSS 16.02fF
C7 XA3/XA5/MP3/a_216_n18# XA3/CN0 0.02fF
C8 XA8/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C9 XDAC1/XC32a<0>/C1A D<6> 0.04fF
C10 XA2/XA5/MP3/a_216_n18# AVDD 0.07fF
C11 XA8/XA4/A XA20/XA3/CO 0.02fF
C12 XA0/CP0 D<7> 2.52fF
C13 XA4/XA1/XA4/MP0/a_216_n18# XA4/XA1/XA2/MP0/a_216_n18# 0.01fF
C14 XA5/XA9/Y XA5/XA9/MN1/S 0.12fF
C15 XA4/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C16 XA4/XA9/B XA4/XA9/MP1/a_216_334# 0.08fF
C17 XA7/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C18 XA5/XA1/XA5/MN2/S XA5/XA1/XA5/MN1/S 0.04fF
C19 XA8/EN XA7/XA1/XA4/MN1/S 0.01fF
C20 D<0> XA8/XA9/A 0.01fF
C21 EN XA0/XA1/XA2/Y 0.21fF
C22 XA4/XA4/A XA4/XA5/MP0/a_216_n18# 0.08fF
C23 XA8/XA9/MN1/a_324_334# XA8/XA11/MN0/a_324_n18# 0.01fF
C24 XA0/XA1/XA1/MP3/a_216_n18# XA0/XA1/XA1/MP2/a_216_n18# 0.01fF
C25 XA3/XA1/XA1/MP2/S XA3/EN 0.01fF
C26 VREF XA8/CN0 0.56fF
C27 XA20/CPO XA20/XA2a/MN1/a_324_n18# 0.01fF
C28 XA1/XA1/XA5/MP2/S XA1/XA2/A 0.06fF
C29 XA1/XA2/MN3/a_324_n18# XA1/CN1 0.03fF
C30 XA4/XA4/MP2/a_216_n18# AVDD 0.07fF
C31 XA3/XA9/MP1/a_216_334# XA3/XA9/B 0.08fF
C32 XA7/XA1/XA4/MN2/S AVSS 0.06fF
C33 XA8/ENO XA8/XA1/XA2/Y 0.10fF
C34 XDAC1/XC32a<0>/XRES16/B D<3> 0.02fF
C35 XA20/XA12/MP0/a_216_n18# XA20/XA12/Y 0.01fF
C36 XA3/XA1/XA4/MN1/S XA3/XA1/XA2/Y 0.05fF
C37 XB1/XA4/MN1/a_324_n18# XB1/XA4/MN0/a_324_n18# 0.01fF
C38 XA20/XA9/Y XA20/XA3/MN0/a_324_n18# 0.08fF
C39 XA20/CPO XA3/CN1 0.21fF
C40 XA6/XA1/XA4/MP2/S AVDD 0.11fF
C41 XB1/XA3/MP0/S XB1/XA3/MN2/a_324_n18# 0.09fF
C42 XA0/XA11/MP1/a_216_n18# XA0/XA11/MP0/a_216_n18# 0.01fF
C43 XDAC1/XC1/XRES1B/B XB1/XA4/GNG 0.03fF
C44 XA8/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C45 XA0/XA1/XA1/MN2/S AVSS 0.30fF
C46 XA7/XA4/A XA20/CNO 0.21fF
C47 XA5/EN XA4/EN 0.06fF
C48 XDAC1/X16ab/XRES8/B SARP 11.94fF
C49 XA8/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C50 XA6/CP0 XA7/EN 0.06fF
C51 XDAC1/XC64b<1>/XRES16/B XDAC1/XC64b<1>/XRES1A/B 1.60fF
C52 XA7/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C53 XA4/XA4/MN3/a_324_n18# XA4/XA4/MN2/a_324_n18# 0.01fF
C54 XA4/XA9/B XA4/CN0 0.07fF
C55 XDAC2/XC32a<0>/XRES4/B XDAC2/XC32a<0>/XRES8/B 2.60fF
C56 XB2/M4/G CK_SAMPLE_BSSW 0.02fF
C57 XA6/XA4/A AVDD 1.42fF
C58 XDAC2/XC64b<1>/XRES4/B XDAC2/XC0/XRES4/B 0.10fF
C59 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC0/XRES8/B 0.02fF
C60 XA8/XA4/MP3/a_216_n18# XA8/XA4/MP2/a_216_n18# 0.01fF
C61 XA3/CN0 D<6> 0.01fF
C62 XA2/XA9/MN0/a_324_n18# XA2/XA9/A 0.15fF
C63 XA20/XA2a/MN2/a_324_n18# XA20/XA2a/MN1/a_324_n18# 0.01fF
C64 XA3/XA1/XA4/MN2/S XA20/CNO 0.01fF
C65 SAR_IN SAR_IP 0.02fF
C66 XA1/XA4/A VREF 0.37fF
C67 D<2> XA20/CPO 0.06fF
C68 XA4/XA1/XA1/MP2/S XA5/EN 0.14fF
C69 XA5/XA2/A XA20/CNO 0.04fF
C70 XA20/XA12/Y XA20/XA10/MP1/a_216_n18# 0.07fF
C71 XA6/XA3/MP2/a_216_n18# VREF 0.03fF
C72 XA1/XA1/XA1/MP3/G XA1/XA1/XA1/MP3/a_216_n18# 0.07fF
C73 XDAC2/XC64a<0>/XRES8/B XDAC2/XC32a<0>/XRES8/B 0.21fF
C74 XA1/XA3/MN0/a_324_n18# XA1/XA3/MN1/a_324_n18# 0.01fF
C75 XA7/CN0 XA20/CPO 0.07fF
C76 XA1/XA9/B XA0/CEO 0.02fF
C77 XA2/CN0 XA5/EN 0.10fF
C78 XA5/CN0 XA4/CN0 4.05fF
C79 XA5/CP0 XA5/CN1 0.03fF
C80 XA0/CP0 VREF 0.83fF
C81 XA3/XA11/MN1/a_324_n18# XA3/XA11/A 0.07fF
C82 XA5/XA4/A XA4/XA4/A 0.03fF
C83 XA5/XA1/XA2/Y XA5/XA1/XA5/MN1/a_324_n18# 0.08fF
C84 XA5/XA6/MP1/S VREF 0.04fF
C85 XA2/XA4/A XA2/XA4/MP0/a_216_n18# 0.07fF
C86 D<3> XA20/CPO 0.07fF
C87 XA5/XA2/MP2/a_216_n18# VREF 0.03fF
C88 XA0/XA8/MP0/a_216_n18# XA1/EN 0.08fF
C89 XA1/XA8/MN0/a_324_n18# XA1/XA7/MN0/a_324_n18# 0.01fF
C90 XDAC2/XC64b<1>/XRES16/B XDAC2/X16ab/XRES1B/B 0.05fF
C91 XA2/XA6/MN3/S AVDD 0.01fF
C92 XA0/XA3/MN0/a_324_n18# XA0/XA2/A 0.07fF
C93 XA6/XA2/A XA5/XA4/A 0.03fF
C94 XA0/XA4/A XA0/XA3/MN2/a_324_n18# 0.01fF
C95 XA6/XA9/A XA6/XA9/MN1/a_324_n18# 0.07fF
C96 XA4/XA1/XA4/MN2/S AVSS 0.06fF
C97 XA0/XA11/A XA0/XA11/MP0/a_216_n18# 0.07fF
C98 XA20/XA9/Y AVDD 2.54fF
C99 XA2/EN XA1/CN0 0.19fF
C100 XB1/XCAPB1/XCAPB2/m3_9828_132# XB1/XA4/GNG 0.04fF
C101 XA20/CNO XA0/CN0 0.05fF
C102 XA4/XA1/XA4/MP0/a_216_n18# XA5/EN 0.08fF
C103 XDAC2/XC128b<2>/XRES4/B XDAC2/XC128b<2>/XRES16/B 0.25fF
C104 XDAC2/XC1/XRES4/B XB2/XA3/B 0.03fF
C105 XA2/CP0 XDAC1/X16ab/XRES16/B 0.03fF
C106 XA1/CEO AVDD 0.75fF
C107 XA7/XA2/MN0/a_324_n18# XA7/EN 0.07fF
C108 XA1/XA1/XA2/Y AVSS 0.27fF
C109 XA8/XA1/XA5/MN1/a_324_n18# XA8/XA1/XA5/MN0/a_324_n18# 0.01fF
C110 D<5> XA3/XA3/MP3/a_216_n18# 0.02fF
C111 XA3/CN0 SARP 0.02fF
C112 XDAC2/XC0/XRES16/B XDAC2/XC0/XRES8/B 1.42fF
C113 XA3/XA1/XA4/MN2/S XA3/XA1/XA4/MN1/S 0.04fF
C114 XDAC1/XC1/XRES8/B XDAC1/XC1/XRES2/B 1.58fF
C115 XDAC2/XC1/XRES4/B AVSS 5.45fF
C116 XA4/XA4/MP1/a_216_n18# XA4/XA4/A 0.15fF
C117 SARN XB1/M6/a_324_n18# 0.02fF
C118 XA8/ENO XA8/CP0 0.06fF
C119 XA4/XA12/A VREF 0.03fF
C120 XA8/XA1/XA5/MN1/a_324_n18# XA20/CNO 0.07fF
C121 XB2/XA4/GNG XB2/M4/G 0.25fF
C122 XA2/XA1/XA1/MP2/S XA2/XA1/XA1/MP3/S 0.04fF
C123 XA0/CP1 XA1/CN1 0.18fF
C124 XA8/XA5/MP0/a_216_n18# VREF 0.02fF
C125 XA7/XA1/XA4/MN2/a_324_n18# XA7/EN 0.08fF
C126 D<1> XA1/CP0 0.04fF
C127 XA0/CEIN XB1/XA1/MP0/G 0.04fF
C128 AVDD XA3/XA5/MP0/a_216_n18# 0.08fF
C129 XDAC1/XC0/XRES4/B SARP 6.32fF
C130 XA6/XA1/XA2/MP0/a_216_n18# XA6/XA1/XA1/MP3/G 0.08fF
C131 XA0/XA6/MN3/S XA0/XA9/B 0.09fF
C132 XA20/XA2a/MP1/a_216_n18# XA20/XA3/CO 0.16fF
C133 XA6/XA1/XA5/MN0/a_324_n18# XA6/EN 0.07fF
C134 EN XA0/XA1/XA1/MN2/S 0.04fF
C135 XA1/XA6/MN3/S AVSS 0.13fF
C136 XA0/XA6/MP1/a_216_n18# AVDD 0.08fF
C137 XA20/XA10/MP1/a_216_n18# CK_SAMPLE 0.01fF
C138 XA4/XA9/MN1/a_324_n18# XA4/XA9/MN0/a_324_n18# 0.01fF
C139 XA3/XA1/XA1/MP0/a_216_n18# XA3/XA1/XA1/MP1/a_216_n18# 0.01fF
C140 XA8/XA11/A XA8/XA9/B 0.03fF
C141 XA20/XA9/A AVDD 1.70fF
C142 XA2/CP0 XA2/XA1/XA1/MP3/G 0.02fF
C143 XA8/ENO XA8/XA9/A 0.08fF
C144 AVDD XA8/XA5/MP3/a_216_n18# 0.08fF
C145 XA8/XA1/XA5/MN1/S AVSS 0.10fF
C146 XA4/XA5/MP1/a_216_n18# XA4/CP0 0.15fF
C147 SARP XB1/XA4/GNG 2.18fF
C148 XA4/XA4/MP0/a_216_n18# XA4/CN1 0.08fF
C149 XDAC1/XC32a<0>/XRES8/B XDAC1/XC128a<1>/XRES1A/B 0.03fF
C150 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC128a<1>/XRES1B/B 0.03fF
C151 XA1/XA1/XA1/MP3/S XA1/XA1/XA1/MP3/G 0.04fF
C152 XA1/XA3/MP0/a_216_n18# XA1/XA2/A 0.08fF
C153 XA8/XA1/XA5/MP1/S EN 0.03fF
C154 XA20/XA3a/A XA20/XA3a/MP0/a_216_n18# 0.08fF
C155 XA0/XA1/XA1/MP3/G AVSS 0.12fF
C156 XA1/XA12/A XA1/XA9/Y 0.02fF
C157 SAR_IN XB2/M4/G 0.65fF
C158 XA2/XA2/MN2/a_324_n18# XA2/CN1 0.02fF
C159 XA2/XA6/MP3/a_216_n18# AVDD 0.08fF
C160 XA6/XA12/A AVDD 0.44fF
C161 XA5/XA4/MN1/a_324_n18# XA5/XA4/MN2/a_324_n18# 0.01fF
C162 XA2/EN XA3/EN 0.06fF
C163 XA5/XA1/XA5/MP1/S XA20/CNO 0.01fF
C164 XA20/XA1/MN4/a_324_n18# XA20/XA1/MN3/a_324_n18# 0.01fF
C165 AVDD XB1/XA5b/MN1/a_324_n18# 0.01fF
C166 XA4/XA4/A VREF 0.37fF
C167 XA8/EN XA20/CPO 0.74fF
C168 XDAC2/XC64b<1>/XRES2/B XDAC2/XC0/XRES2/B 0.05fF
C169 XA8/CN0 XA8/CP0 0.46fF
C170 XA4/XA5/MN3/a_324_n18# XA4/CN0 0.01fF
C171 XA7/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C172 XB2/CKN XB2/XA3/MP0/a_216_334# 0.09fF
C173 D<5> AVDD 1.85fF
C174 XA2/XA4/MP1/a_216_n18# XA2/XA4/MP2/a_216_n18# 0.01fF
C175 XA1/XA1/XA1/MP2/a_216_n18# XA20/CPO 0.06fF
C176 XDAC1/XC128a<1>/XRES2/B XDAC1/XC128a<1>/XRES4/B 0.55fF
C177 XA6/XA2/A VREF 0.36fF
C178 XA4/XA11/A VREF 0.02fF
C179 XA0/CEO XA0/XA11/MP1/S 0.02fF
C180 D<7> XA1/XA3/MN3/a_324_n18# 0.02fF
C181 XB1/XA4/MP1/a_216_n18# XB1/XA4/MP1/a_216_334# 0.01fF
C182 XA0/XA9/B XA0/XA11/A 0.03fF
C183 D<8> AVSS 3.59fF
C184 XA5/XA3/MN2/a_324_n18# XA5/XA4/A 0.01fF
C185 XB2/XA5b/MN1/a_324_n18# CK_SAMPLE_BSSW 0.01fF
C186 XA3/XA1/XA4/MP1/S AVDD 0.14fF
C187 XA2/CN1 XA2/XA2/MN1/a_324_n18# 0.03fF
C188 XB1/XA7/MP1/a_216_334# XB1/XA7/MP1/a_216_n18# 0.01fF
C189 XDAC1/XC64a<0>/XRES1B/B XDAC1/XC64a<0>/XRES1A/B 0.01fF
C190 XA6/XA5/MP0/a_216_n18# XA6/XA4/A 0.08fF
C191 XA4/XA1/XA1/MN1/a_324_n18# XA4/EN 0.08fF
C192 XA1/CP0 XA3/CN1 0.13fF
C193 SARN XDAC2/XC32a<0>/XRES16/B 21.65fF
C194 XA8/EN XA8/XA1/XA4/MN2/S 0.02fF
C195 XA1/CP0 XA1/XA5/MP2/a_216_n18# 0.15fF
C196 XA3/XA1/XA1/MN2/S AVDD 0.05fF
C197 XA6/XA1/XA1/MN0/a_324_n18# AVSS 0.08fF
C198 XA2/EN XA2/XA1/XA1/MN2/S 0.05fF
C199 VREF CK_SAMPLE_BSSW 0.03fF
C200 XA3/XA12/MP0/a_216_n18# XA2/CEO 0.08fF
C201 XDAC2/X16ab/XRES1B/B SARN 1.79fF
C202 XA2/XA4/A AVSS 1.07fF
C203 XDAC1/XC64b<1>/XRES16/B XDAC1/XC64b<1>/XRES2/B 1.61fF
C204 XA1/XA1/XA2/Y EN 0.07fF
C205 XA1/XA1/XA5/MP1/S EN 0.03fF
C206 XA5/XA7/MP0/a_216_n18# XA5/XA6/MP3/a_216_n18# 0.01fF
C207 XDAC2/XC128a<1>/XRES4/B XDAC2/XC32a<0>/XRES4/B 0.10fF
C208 XA4/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C209 XA7/XA1/XA2/Y XA8/XA1/XA2/Y 0.02fF
C210 AVDD XA2/XA1/XA5/MP0/a_216_n18# 0.08fF
C211 XA20/XA3/MN6/a_324_n18# XA20/XA3/N2 0.01fF
C212 XA4/CP0 AVDD 1.31fF
C213 XA3/XA9/A XA3/XA9/MP1/a_216_n18# 0.08fF
C214 D<2> XA1/CP0 0.05fF
C215 XA1/XA6/MN3/S CK_SAMPLE 0.03fF
C216 XA1/XA1/XA1/MN0/a_324_n18# XA1/XA1/XA1/MN1/a_324_n18# 0.01fF
C217 XA8/XA11/A VREF 0.02fF
C218 XA3/XA1/XA5/MN2/S AVDD 0.02fF
C219 D<6> XA20/CNO 0.05fF
C220 XA8/XA1/XA1/MP1/a_216_n18# XA8/XA1/XA1/MP3/G 0.01fF
C221 XA7/CP0 AVSS 0.91fF
C222 XA0/XA4/A XA20/CNO 0.17fF
C223 XA3/XA12/A VREF 0.03fF
C224 XDAC2/XC0/XRES1B/B XDAC2/XC0/XRES8/B 0.12fF
C225 XA20/XA3/MN6/a_324_n18# XA20/XA4/MN0/a_324_n18# 0.01fF
C226 XA20/XA9/Y XA20/XA3/MP2/a_216_n18# 0.08fF
C227 XA20/XA9/MP0/a_216_334# XA20/XA11/Y 0.06fF
C228 XB1/M4/G XB1/XA4/MP1/a_216_334# 0.08fF
C229 XA7/XA1/XA2/Y XA7/XA1/XA5/MN0/a_324_n18# 0.02fF
C230 XA6/XA3/MP0/a_216_n18# XA6/XA2/MP3/a_216_n18# 0.01fF
C231 XA1/CP0 D<3> 0.04fF
C232 XA1/XA9/MP1/a_216_334# XA1/XA9/Y 0.07fF
C233 XDAC1/XC1/XRES4/B XDAC1/XC64a<0>/XRES1A/B 0.01fF
C234 XA3/XA2/MP3/a_216_n18# VREF 0.03fF
C235 XA8/XA1/XA5/MN1/S EN 0.01fF
C236 XA6/XA6/MP0/a_216_n18# AVDD 0.08fF
C237 XA7/XA2/MN2/a_324_n18# XA7/XA2/MN1/a_324_n18# 0.01fF
C238 XA4/CN1 AVSS 0.79fF
C239 XA6/EN XA5/XA1/XA1/MP3/S 0.10fF
C240 XA8/EN XA7/XA8/MP0/a_216_n18# 0.08fF
C241 EN XA0/XA1/XA1/MP3/G 0.13fF
C242 XA6/EN XA5/XA1/XA1/MN2/a_324_n18# 0.01fF
C243 XA4/EN XA3/XA1/XA1/MN1/a_324_n18# 0.01fF
C244 XDAC2/XC64b<1>/XRES16/B XA1/CN1 0.17fF
C245 XA3/XA9/B XA4/EN 0.07fF
C246 XA3/CN0 XDAC2/X16ab/XRES16/B 0.02fF
C247 XB1/M4/G XB1/XA4/MP1/a_216_n18# 0.08fF
C248 XA3/DONE AVSS 0.15fF
C249 D<1> XA7/XA6/MP1/a_216_n18# 0.01fF
C250 XA6/EN AVSS 1.54fF
C251 XA3/XA8/MN0/a_324_n18# XA3/XA9/B 0.01fF
C252 XA8/XA4/MP0/a_216_n18# XA8/XA4/A 0.07fF
C253 XA8/XA1/XA4/MP2/S EN 0.02fF
C254 XB2/XA5/MN1/a_324_334# AVSS 0.10fF
C255 XB2/XA4/GNG XB2/XA1/MP0/G 0.06fF
C256 XA20/XA2/MP4/a_216_n18# XA20/XA3a/A 0.01fF
C257 XB2/M2/a_324_n18# SAR_IN 0.02fF
C258 XA8/XA5/MP0/a_216_n18# XA8/CP0 0.07fF
C259 XA20/XA4/MP0/S XA20/XA4/MN6/a_324_n18# 0.01fF
C260 AVDD XB1/XA4/MP1/a_216_334# 0.09fF
C261 XA3/CN0 XA4/CN0 2.51fF
C262 XA5/XA12/A AVSS 0.39fF
C263 EN D<8> 0.30fF
C264 D<4> XA3/CP0 1.94fF
C265 XA8/EN XA7/XA1/XA2/MN0/a_324_n18# 0.09fF
C266 XA8/XA1/XA5/MP2/S AVDD 0.08fF
C267 XDAC2/XC1/XRES1A/B SARN 1.51fF
C268 XA6/CN0 XA6/CN1 0.08fF
C269 XA0/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C270 XA6/XA1/XA4/MP1/S XA20/CPO 0.02fF
C271 XA6/XA11/MN0/a_324_n18# AVSS 0.01fF
C272 XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MP3/S 0.04fF
C273 XA6/EN XA5/XA9/B 0.07fF
C274 XA3/CN0 XA5/CN0 0.14fF
C275 XA20/XA3/MP6/a_216_n18# XA20/XA3/CO 0.01fF
C276 XA1/XA3/MP0/a_216_n18# XA1/CN1 0.07fF
C277 D<1> XA7/XA9/A 0.01fF
C278 XA8/XA4/MN2/a_324_n18# XA8/CP0 0.01fF
C279 XA2/XA4/A EN 0.10fF
C280 XA3/XA2/A XA4/XA4/A 0.03fF
C281 XA1/XA4/MN3/a_324_n18# XA1/XA4/MN2/a_324_n18# 0.01fF
C282 XA7/DONE XA7/XA9/Y 0.06fF
C283 XA1/XA1/XA1/MP3/G XA20/CPO 0.15fF
C284 XA7/CP0 CK_SAMPLE 0.09fF
C285 AVDD XB1/XA4/MP1/a_216_n18# 0.09fF
C286 XA0/XA5/MP0/a_216_n18# VREF 0.02fF
C287 XA2/XA4/MN3/a_324_n18# XA2/XA4/A 0.15fF
C288 XA5/XA9/B XA5/XA12/A 0.01fF
C289 XDAC1/XC128a<1>/XRES1B/B XDAC1/XC128b<2>/XRES16/B 0.05fF
C290 SAR_IN XB2/XA1/MP0/G 0.01fF
C291 XA8/XA2/MP3/a_216_n18# XA8/XA3/MP0/a_216_n18# 0.01fF
C292 XA8/XA7/MN0/a_324_n18# XA8/XA6/MN3/a_324_n18# 0.01fF
C293 XDAC2/XC1/XRES1B/B XDAC2/XC1/XRES1A/B 0.01fF
C294 XA0/XA9/A AVDD 0.62fF
C295 XA2/XA2/MP2/a_216_n18# AVDD 0.07fF
C296 XDAC1/XC64a<0>/XRES4/B SARP 6.32fF
C297 XA2/CP0 XA3/CP0 0.97fF
C298 XA4/XA6/MP1/a_216_n18# XA4/XA6/MP0/a_216_n18# 0.01fF
C299 XA6/XA6/MP1/S VREF 0.04fF
C300 XA1/XA1/XA1/MP2/S XA1/EN 0.01fF
C301 XA0/XA1/XA5/MN2/S AVSS 0.09fF
C302 D<3> XA5/XA6/MP2/a_216_n18# 0.07fF
C303 XA3/EN XA2/XA1/XA1/MN3/a_324_n18# 0.01fF
C304 AVDD XA2/XA1/XA5/MP2/a_216_n18# 0.08fF
C305 XA2/CN0 XA1/CN1 0.08fF
C306 XA7/EN XA20/CNO 0.93fF
C307 XA3/EN XA2/XA1/XA2/MP0/a_216_n18# 0.08fF
C308 XA4/XA11/MP0/a_216_n18# XA4/XA9/MP1/a_216_334# 0.01fF
C309 XA3/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C310 XA8/XA11/MP1/a_216_n18# XA7/CEO 0.06fF
C311 XA3/XA5/MP2/a_216_n18# XA3/CP0 0.15fF
C312 XA4/XA5/MP1/a_216_n18# AVDD 0.07fF
C313 XA3/XA3/MP3/a_216_n18# AVDD 0.07fF
C314 XA5/XA9/Y XA5/XA9/A 0.04fF
C315 XA7/EN XA6/XA1/XA1/MP3/S 0.10fF
C316 XA1/XA6/MP1/a_216_n18# XA1/XA6/MP2/a_216_n18# 0.01fF
C317 XA3/XA11/A XA3/XA11/MN0/a_324_n18# 0.09fF
C318 XA4/EN XA3/XA1/XA1/MN3/a_324_n18# 0.02fF
C319 XA8/XA3/MP2/a_216_n18# XA8/CN1 0.15fF
C320 XA7/XA2/MP3/a_216_n18# XA7/XA3/MP0/a_216_n18# 0.01fF
C321 XA8/XA7/MN0/a_324_n18# XA8/XA9/B 0.01fF
C322 XA6/XA9/Y XA6/XA11/MN0/a_324_n18# 0.07fF
C323 XA3/XA1/XA4/MP0/a_216_n18# XA3/XA1/XA4/MP1/a_216_n18# 0.01fF
C324 XA7/XA12/A XA7/CEO 0.21fF
C325 XA4/CP0 XA5/EN 0.06fF
C326 XA6/EN CK_SAMPLE 0.09fF
C327 XA8/XA5/MN3/a_324_n18# XA8/CP0 0.15fF
C328 XA20/XA9/MN0/a_324_n18# XA20/XA4/MN6/a_324_n18# 0.01fF
C329 D<1> XA7/XA1/XA1/MP3/G 0.02fF
C330 SARN XB1/XA1/Y 0.03fF
C331 XA1/XA9/MP1/a_216_n18# XA1/XA9/MP0/a_216_n18# 0.01fF
C332 XA4/CN1 EN 0.05fF
C333 XA4/XA13/MN1/a_324_n18# XA4/XA12/A 0.07fF
C334 XA0/XA5/MP1/a_216_n18# AVDD 0.07fF
C335 EN XA2/XA1/XA4/MP1/a_216_n18# 0.15fF
C336 AVDD XA2/XA1/XA4/MP0/a_216_n18# 0.08fF
C337 XA0/CP1 AVSS 3.39fF
C338 SARN XB1/CKN 0.01fF
C339 XA2/XA6/MP3/S XA3/EN 0.02fF
C340 XA1/XA2/MN2/a_324_n18# XA1/XA2/MN1/a_324_n18# 0.01fF
C341 XA7/XA4/MN0/a_324_n18# XA7/CN1 0.07fF
C342 XDAC2/XC128b<2>/XRES8/B XDAC2/X16ab/XRES1A/B 0.03fF
C343 XDAC2/XC128b<2>/XRES1B/B XDAC2/X16ab/XRES1B/B 0.03fF
C344 XDAC2/XC64b<1>/XRES1A/B XDAC2/XC64b<1>/XRES1B/B 0.01fF
C345 D<0> XA8/XA7/MP0/a_216_n18# 0.08fF
C346 XA20/XA12/Y XA20/XA11/Y 0.17fF
C347 XA20/XA11/Y AVSS 0.41fF
C348 XB2/XA7/MP1/a_216_n18# XB2/XA4/MP1/a_216_334# 0.01fF
C349 AVDD XB1/M4/G 0.65fF
C350 XA5/XA9/A XA5/XA11/A 0.01fF
C351 SARN XA1/CN1 0.34fF
C352 XA7/CN0 XA7/XA6/MP1/a_216_n18# 0.15fF
C353 XA6/EN EN 1.01fF
C354 XA5/CP0 XA5/CN0 0.60fF
C355 XA5/XA1/XA4/MN2/S XA5/XA1/XA2/Y 0.05fF
C356 XA5/CN0 XA5/XA6/MP1/a_216_n18# 0.15fF
C357 XA8/ENO XA20/CPO 0.37fF
C358 XDAC2/XC128a<1>/XRES16/B XDAC2/XC32a<0>/XRES1B/B 0.05fF
C359 XA1/XA9/MP1/a_216_334# XA1/XA9/MP1/a_216_n18# 0.01fF
C360 EN XA0/XA2/MP0/a_216_n18# 0.08fF
C361 XA6/XA9/MP1/a_216_334# AVDD 0.09fF
C362 XA4/XA2/A XA4/XA4/A 0.14fF
C363 XDAC1/XC64b<1>/XRES16/B XDAC1/X16ab/XRES4/B 0.03fF
C364 XA4/EN XA3/XA1/XA1/MP3/G 0.26fF
C365 D<6> XA2/XA1/XA2/Y 0.02fF
C366 XA1/XA4/A XA1/XA1/XA4/MN1/S 0.02fF
C367 XA20/XA13/MN1/a_324_n18# AVSS 0.09fF
C368 XA3/XA9/A XA3/XA9/MP0/a_216_n18# 0.14fF
C369 XA3/XA2/A XA3/XA2/MP3/a_216_n18# 0.15fF
C370 XA6/XA4/MP0/a_216_n18# XA6/XA4/A 0.07fF
C371 XA6/XA2/MP2/a_216_n18# AVDD 0.07fF
C372 EN XA0/XA1/XA1/MN0/a_324_n18# 0.08fF
C373 XA20/XA2/MN6/a_324_334# XA20/XA3/CO 0.14fF
C374 XA4/XA9/B XA4/XA9/MN1/a_324_334# 0.07fF
C375 XDAC2/XC0/XRES4/B SARP 0.02fF
C376 XA6/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C377 XA4/CP0 XA4/XA5/MN0/a_324_n18# 0.09fF
C378 XA7/XA4/A XA8/XA4/A 0.16fF
C379 XA8/ENO XA20/XA3/N1 0.01fF
C380 XA4/XA13/MN1/a_324_n18# XA4/XA12/MN0/a_324_n18# 0.01fF
C381 XA7/CN0 XA7/XA5/MN1/a_324_n18# 0.02fF
C382 XA5/XA1/XA1/MN2/a_324_n18# XA5/XA1/XA1/MN3/a_324_n18# 0.01fF
C383 XA3/EN XA2/XA1/XA1/MP3/G 0.28fF
C384 XB1/XA3/MP2/a_216_n18# XB1/XA4/MP0/a_216_n18# 0.01fF
C385 XA7/XA1/XA2/Y XA7/XA1/XA4/MN1/S 0.05fF
C386 XDAC1/XC128b<2>/XRES2/B XDAC1/X16ab/XRES2/B 0.05fF
C387 XA6/EN XA5/XA1/XA2/MN0/a_324_n18# 0.09fF
C388 XA8/XA11/A XA8/XA9/A 0.01fF
C389 XA5/XA1/XA5/MN2/a_324_n18# XA5/XA1/XA5/MN1/a_324_n18# 0.01fF
C390 XA3/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C391 XA0/CP0 XDAC1/XC64b<1>/XRES16/B 0.02fF
C392 XA6/XA3/MP3/a_216_n18# VREF 0.03fF
C393 XA7/XA1/XA1/MP0/a_216_n18# AVDD 0.14fF
C394 XA2/CN0 XA3/XA1/XA1/MP3/G 0.01fF
C395 XA6/XA6/MP1/a_216_n18# XA6/XA6/MP2/a_216_n18# 0.01fF
C396 XA7/XA12/A XA7/XA9/B 0.01fF
C397 XA5/XA3/MP1/a_216_n18# XA5/CN1 0.15fF
C398 XA0/XA9/A XA0/XA8/MN0/a_324_n18# 0.09fF
C399 XA0/XA2/MP1/a_216_n18# AVDD 0.08fF
C400 SARP XB1/XA3/MP0/S 0.02fF
C401 XA1/XA1/XA5/MN2/S AVDD 0.02fF
C402 XA5/XA2/A XA5/XA1/XA5/MN2/S 0.05fF
C403 XA2/EN XA1/XA1/XA4/MP0/a_216_n18# 0.08fF
C404 XA6/CN0 XA1/CN0 0.20fF
C405 XDAC1/XC32a<0>/XRES16/B XA0/CP0 0.05fF
C406 XA3/XA9/Y AVDD 0.58fF
C407 XA0/XA1/XA5/MN0/a_324_n18# XA0/XA1/XA2/Y 0.02fF
C408 EN XA0/XA1/XA5/MN2/S 0.02fF
C409 XA2/CP0 XA2/XA6/MN0/a_324_n18# 0.07fF
C410 XB2/XCAPB1/XCAPB1/m3_252_308# XB2/XA3/B 0.02fF
C411 XA20/CPO XA2/XA1/XA1/MN2/a_324_n18# 0.08fF
C412 XA6/XA5/MN1/a_324_n18# XA6/CP0 0.15fF
C413 XA20/CPO XA2/XA1/XA4/MP1/S 0.02fF
C414 EN XA5/XA1/XA5/MP2/a_216_n18# 0.16fF
C415 XA4/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C416 XA4/XA1/XA2/Y AVDD 0.33fF
C417 XA5/XA11/MN1/a_324_n18# XA4/CEO 0.08fF
C418 XA4/XA13/MP1/a_216_334# AVDD 0.17fF
C419 XA2/XA1/XA5/MN2/S AVSS 0.09fF
C420 XA6/XA6/MN2/a_324_n18# XA6/XA6/MN3/a_324_n18# 0.01fF
C421 XA2/XA1/XA1/MN2/S XA2/XA1/XA1/MP3/G 0.08fF
C422 XA2/XA13/MN1/a_324_n18# AVSS 0.09fF
C423 XA0/CP1 CK_SAMPLE 0.10fF
C424 XA4/XA1/XA1/MP2/a_216_n18# XA20/CPO 0.06fF
C425 XA0/XA1/XA4/MN1/S AVSS 0.10fF
C426 XA3/XA6/MP0/a_216_n18# VREF 0.01fF
C427 XDAC2/XC1/XRES8/B XDAC2/XC64a<0>/XRES16/B 0.03fF
C428 XA6/XA6/MP3/a_216_n18# AVDD 0.08fF
C429 XA6/XA4/MP1/a_216_n18# VREF 0.02fF
C430 XA20/XA11/Y CK_SAMPLE 0.08fF
C431 XA4/XA9/MN1/S AVDD 0.01fF
C432 XA2/XA4/A XA2/XA4/MP3/a_216_n18# 0.15fF
C433 XA8/XA2/A XA20/XA3/CO 0.05fF
C434 XA7/XA8/MP0/a_216_n18# XA7/XA7/MP0/a_216_n18# 0.01fF
C435 XA7/XA6/MN2/a_324_n18# XA7/XA6/MN3/a_324_n18# 0.01fF
C436 XA8/XA1/XA4/MP0/a_216_n18# XA8/XA1/XA2/MP0/a_216_n18# 0.01fF
C437 XA7/XA1/XA1/MP3/G XA7/CN0 0.02fF
C438 XA1/XA9/MN1/S AVDD 0.01fF
C439 XA4/CN0 XA20/CNO 0.06fF
C440 XA7/XA11/A AVDD 0.45fF
C441 XA2/XA3/MP1/a_216_n18# D<6> 0.02fF
C442 XA6/CP0 XA5/CP0 0.03fF
C443 XA5/XA7/MN0/a_324_n18# AVSS 0.01fF
C444 XA1/XA1/XA2/Y XA2/CN1 0.03fF
C445 XA1/XA9/A XA0/XA9/A 0.01fF
C446 XA0/CP1 EN 0.08fF
C447 XA8/XA1/XA1/MP3/G XA8/XA1/XA2/MP0/a_216_n18# 0.08fF
C448 XA1/XA4/A XA20/CPO 0.03fF
C449 XA1/CP0 XA1/XA1/XA1/MP3/G 0.02fF
C450 XB1/XA3/MP0/a_216_n18# XB1/XA0/MP0/a_216_n18# 0.01fF
C451 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC0/XRES16/B 0.05fF
C452 XA3/EN XA3/XA4/A 0.20fF
C453 XA5/CN0 XA20/CNO 0.06fF
C454 XA0/XA1/XA2/MN0/a_324_n18# XA0/XA1/XA1/MN3/a_324_n18# 0.01fF
C455 XA5/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C456 XA7/XA5/MN2/a_324_n18# XA7/XA5/MN3/a_324_n18# 0.01fF
C457 XA20/XA1/MP0/S SARP 0.21fF
C458 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC64a<0>/XRES2/B 0.23fF
C459 XA5/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C460 XA6/XA9/A XA7/EN 0.09fF
C461 XA2/XA6/MP1/a_216_n18# XA2/XA6/MP2/a_216_n18# 0.01fF
C462 XA2/XA8/MP0/a_216_n18# XA2/XA9/MP0/a_216_n18# 0.01fF
C463 XB2/CKN XB2/XA4/MP1/a_216_n18# 0.08fF
C464 XA5/XA7/MN0/a_324_n18# XA5/XA9/B 0.01fF
C465 XA0/CP0 XA20/CPO 0.05fF
C466 XA8/XA1/XA1/MP3/a_216_n18# AVDD 0.09fF
C467 XA7/XA2/MP2/a_216_n18# XA7/XA2/MP3/a_216_n18# 0.01fF
C468 XA5/XA5/MP1/a_216_n18# XA5/XA5/MP0/a_216_n18# 0.01fF
C469 XA5/XA2/MN3/a_324_n18# XA5/XA2/MN2/a_324_n18# 0.01fF
C470 XA0/XA2/MN0/a_324_n18# XA0/XA2/MN1/a_324_n18# 0.01fF
C471 XA7/XA1/XA1/MN2/S XA7/XA1/XA1/MP3/G 0.08fF
C472 XDAC2/XC64b<1>/XRES16/B AVSS 16.03fF
C473 AVDD XA20/XA4/MP3_DMY/a_216_n18# 0.24fF
C474 XB2/XA3/B XB2/XA3/MP0/a_216_n18# 0.01fF
C475 XA6/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C476 XA0/XA6/MN2/a_324_n18# XA0/XA6/MN3/a_324_n18# 0.01fF
C477 XA8/EN XA7/XA9/A 0.09fF
C478 XA4/XA12/MP0/a_216_n18# AVDD 0.08fF
C479 XA1/XA1/XA5/MP2/S EN 0.04fF
C480 XA2/XA3/MN0/a_324_n18# XA2/CN1 0.10fF
C481 XA1/XA6/MP0/a_216_n18# XA1/CN0 0.08fF
C482 XA0/XA3/MP1/a_216_n18# VREF 0.02fF
C483 XA7/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C484 XDAC2/XC64a<0>/XRES1A/B XDAC2/XC64a<0>/XRES8/B 0.12fF
C485 XA7/XA3/MP2/a_216_n18# XA7/XA3/MP1/a_216_n18# 0.01fF
C486 XB2/XCAPB1/XCAPB4/m3_324_308# XB2/XA3/B 0.02fF
C487 XDAC1/XC1/XRES4/B XB1/XA3/B 0.03fF
C488 XA8/ENO XA8/XA7/MP0/a_216_n18# 0.07fF
C489 XA5/XA1/XA4/MN2/S XA5/XA1/XA4/MN1/S 0.04fF
C490 XA5/XA2/A XA5/XA1/XA5/MP2/S 0.06fF
C491 XA6/XA12/MP0/a_216_n18# XA6/XA11/MP1/a_216_n18# 0.01fF
C492 XA0/XA9/MP1/a_216_n18# XA0/XA9/MP1/a_216_334# 0.01fF
C493 XA5/XA11/MP0/a_216_n18# AVDD 0.09fF
C494 XA3/CP0 XA1/CN0 0.01fF
C495 XA0/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C496 XA7/XA12/A AVSS 0.39fF
C497 AVDD XA6/XA1/XA1/MP3/a_216_n18# 0.08fF
C498 D<5> XA3/XA9/B 0.05fF
C499 XDAC1/XC128a<1>/XRES1B/B XDAC1/XC128b<2>/XRES1B/B 0.03fF
C500 XA4/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C501 XA8/XA11/MN1/a_324_n18# XA8/XA11/A 0.07fF
C502 XA8/XA9/MN1/a_324_334# XA8/XA9/B 0.07fF
C503 XB1/XCAPB1/XCAPB3/m3_324_308# XB1/XA4/GNG 0.07fF
C504 XA20/XA3/MP2/a_216_n18# AVDD 0.15fF
C505 XA5/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C506 XA5/EN AVDD 4.84fF
C507 XA2/CN1 D<8> 0.76fF
C508 XA6/XA9/B D<2> 0.05fF
C509 EN XA2/XA1/XA5/MN2/S 0.02fF
C510 XA1/XA1/XA2/Y D<7> 0.02fF
C511 XA20/XA3/MP5/a_216_n18# AVDD 0.10fF
C512 XA4/EN AVSS 1.44fF
C513 XA8/EN XA7/XA1/XA4/MP0/a_216_n18# 0.08fF
C514 XDAC1/XC0/XRES1B/B XDAC1/XC0/XRES8/B 0.12fF
C515 EN XA0/XA1/XA4/MN1/S 0.02fF
C516 XA5/XA1/XA1/MN3/a_324_n18# XA5/XA1/XA2/MN0/a_324_n18# 0.01fF
C517 XB2/XA2/MP0/G XB2/XA4/GNG 0.07fF
C518 EN XA2/XA2/MP0/a_216_n18# 0.08fF
C519 XA6/XA5/MP0/a_216_n18# AVDD 0.08fF
C520 XA3/XA13/MN1/a_324_n18# XA3/XA12/MN0/a_324_n18# 0.01fF
C521 XA4/XA1/XA1/MP1/a_216_n18# XA4/XA1/XA1/MP2/a_216_n18# 0.01fF
C522 XA1/XA9/A AVDD 0.62fF
C523 XA8/EN XA7/XA1/XA1/MP3/G 0.26fF
C524 XB2/XA3/B XB2/XCAPB1/XCAPB1/m3_324_308# 0.02fF
C525 XA2/XA4/A XA2/CN1 0.62fF
C526 XA6/XA2/A XA6/XA2/MP3/a_216_n18# 0.15fF
C527 XA20/XA2/MP6/a_216_n18# XA20/XA3a/A 0.01fF
C528 XA7/XA1/XA2/Y XA20/CPO 0.24fF
C529 XA3/XA4/MN0/a_324_n18# XA3/XA4/MN1/a_324_n18# 0.01fF
C530 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC128a<1>/XRES8/B 0.02fF
C531 XA7/DONE XA7/XA9/A 0.07fF
C532 XA6/XA3/MN2/a_324_n18# XA6/XA3/MN3/a_324_n18# 0.01fF
C533 XA6/XA1/XA5/MP2/a_216_n18# XA6/XA2/MP0/a_216_n18# 0.01fF
C534 XA5/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C535 XA0/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C536 XA2/EN XA1/XA1/XA4/MN2/S 0.01fF
C537 XA8/XA1/XA5/MP1/S VREF 0.02fF
C538 XA5/EN XA4/XA1/XA2/MP0/a_216_n18# 0.08fF
C539 XA4/XA1/XA2/Y XA5/EN 0.10fF
C540 XA8/XA4/MN2/a_324_n18# XA8/XA4/MN3/a_324_n18# 0.01fF
C541 XA8/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C542 D<5> XA1/CN1 0.04fF
C543 XA6/EN XA6/XA1/XA1/MP3/G 0.03fF
C544 XA4/XA4/A XA20/CPO 0.03fF
C545 XA2/CN0 AVSS 1.01fF
C546 XA2/XA13/MN1/a_324_n18# XA2/XA12/A 0.07fF
C547 XA6/CEO XA6/XA11/MP1/S 0.02fF
C548 XA3/CP0 XA3/EN 0.10fF
C549 XA2/DONE XA2/XA9/A 0.07fF
C550 XA20/XA2/N2 XA20/XA2/MP2/a_216_n18# 0.01fF
C551 XB2/CKN CK_SAMPLE_BSSW 0.12fF
C552 SARP XB1/M8/a_324_n18# 0.01fF
C553 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128a<1>/XRES1B/B 0.12fF
C554 XA3/XA4/MN1/a_324_n18# XA3/XA4/A 0.15fF
C555 XA8/XA1/XA2/Y XA8/XA1/XA4/MN2/a_324_n18# 0.08fF
C556 XA7/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C557 XB2/XA3/B SARN 0.41fF
C558 XA2/XA2/MP1/a_216_n18# XA2/XA2/MP0/a_216_n18# 0.01fF
C559 D<5> XA3/XA6/MP1/a_216_n18# 0.01fF
C560 XA2/CN0 XA2/XA9/B 0.07fF
C561 XA7/XA1/XA5/MP1/S XA7/XA1/XA5/MN1/S 0.01fF
C562 SARN AVSS 113.21fF
C563 XB2/M5/a_324_n18# SARN 0.02fF
C564 AVDD XA7/XA2/A 1.07fF
C565 XDAC2/XC128b<2>/XRES4/B XDAC2/X16ab/XRES16/B 0.03fF
C566 XA1/XA1/XA4/MP1/S XA1/XA1/XA4/MP2/S 0.04fF
C567 XA5/XA1/XA5/MP2/S XA5/XA1/XA5/MP1/S 0.04fF
C568 XA5/XA6/MN1/S AVSS 0.15fF
C569 XDAC2/XC64b<1>/XRES4/B XDAC2/X16ab/XRES4/B 0.10fF
C570 XA8/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C571 XDAC2/XC32a<0>/XRES2/B XDAC2/XC32a<0>/XRES16/B 1.61fF
C572 XA2/XA1/XA4/MN1/S AVSS 0.10fF
C573 XA0/XA9/A XA0/XA9/MP0/a_216_n18# 0.14fF
C574 XA0/XA3/MP0/a_216_n18# XA0/XA3/MP1/a_216_n18# 0.01fF
C575 XDAC1/XC128a<1>/XRES1A/B SARP 1.50fF
C576 D<6> XA2/XA9/A 0.01fF
C577 XA0/XA6/MP0/a_216_n18# VREF 0.01fF
C578 D<7> D<8> 0.05fF
C579 XA0/XA2/MN3/a_324_n18# XA0/XA3/MN0/a_324_n18# 0.01fF
C580 XDAC1/XC64a<0>/XRES16/B XDAC1/XC64a<0>/XRES1A/B 1.60fF
C581 XDAC2/XC128a<1>/XRES1B/B SARN 1.79fF
C582 XA1/XA1/XA5/MP1/S VREF 0.02fF
C583 XA4/EN CK_SAMPLE 0.08fF
C584 XA7/XA1/XA2/MN0/a_324_n18# XA7/XA1/XA1/MN3/a_324_n18# 0.01fF
C585 XA1/CP0 XA1/XA4/A 0.57fF
C586 XA5/XA5/MP2/a_216_n18# XA5/XA5/MP1/a_216_n18# 0.01fF
C587 CK_SAMPLE XA8/XA6/MN1/a_324_n18# 0.16fF
C588 XDAC2/XC1/XRES1B/B AVSS 2.94fF
C589 XB2/XA5b/MP1/a_216_n18# AVDD 0.16fF
C590 XA4/XA3/MN1/a_324_n18# D<4> 0.02fF
C591 XDAC1/XC128a<1>/XRES16/B XDAC1/XC128b<2>/XRES1A/B 0.04fF
C592 XA8/XA5/MP3/a_216_n18# XA8/XA6/MP0/a_216_n18# 0.01fF
C593 XA5/XA9/B XA5/XA6/MN1/S 0.05fF
C594 EN XA0/XA1/XA4/MP1/a_216_n18# 0.15fF
C595 XA4/EN EN 1.00fF
C596 XA20/CPO XA2/XA1/XA1/MP3/a_216_n18# 0.08fF
C597 XA8/XA11/MP1/a_216_n18# XA8/XA12/MP0/a_216_n18# 0.01fF
C598 D<5> XA3/XA1/XA1/MP3/G 0.02fF
C599 XA1/CP0 XA0/CP0 1.65fF
C600 XA2/XA3/MP0/a_216_n18# AVDD 0.08fF
C601 XA1/XA9/B XA1/XA9/MN1/a_324_n18# 0.09fF
C602 XA2/XA1/XA1/MP2/a_216_n18# XA2/XA1/XA1/MP3/G 0.01fF
C603 XA3/XA13/MN1/a_324_334# AVSS 0.10fF
C604 XA2/CN0 CK_SAMPLE 0.07fF
C605 XDAC2/XC64b<1>/XRES16/B XDAC2/XC0/XRES1A/B 0.04fF
C606 XA20/XA9/A XA20/XA9/MP0/a_216_334# 0.08fF
C607 XA3/XA7/MN0/a_324_n18# XA4/EN 0.08fF
C608 XA3/XA6/MN1/a_324_n18# XA3/XA6/MN2/a_324_n18# 0.01fF
C609 XDAC2/XC64b<1>/XRES8/B XDAC2/XC64b<1>/XRES16/B 1.42fF
C610 XDAC1/XC1/XRES8/B AVSS 9.01fF
C611 XA20/XA3/MN1/a_324_n18# SARN 0.08fF
C612 XA7/XA2/MP0/a_216_n18# XA7/XA1/XA5/MP2/a_216_n18# 0.01fF
C613 XB2/CKN XB2/XA4/GNG 0.25fF
C614 XA1/XA2/A AVDD 1.07fF
C615 XA20/XA3a/A XA20/XA4/MP0/a_216_n18# 0.08fF
C616 XA3/XA1/XA1/MN0/a_324_n18# XA3/EN 0.09fF
C617 XA5/XA1/XA1/MP3/G XA6/EN 0.26fF
C618 XA2/CP0 XA2/XA2/A 0.04fF
C619 XA1/CEO XA2/XA11/A 0.08fF
C620 XA3/XA8/MN0/a_324_n18# XA3/XA7/MN0/a_324_n18# 0.01fF
C621 XA20/XA11/MN0/a_324_n18# XA20/XA10/MN1/a_324_n18# 0.01fF
C622 XA5/XA1/XA4/MN0/a_324_n18# XA5/XA1/XA2/MN0/a_324_n18# 0.01fF
C623 XDAC1/XC128b<2>/XRES16/B XDAC1/XC128b<2>/XRES1B/B 0.12fF
C624 XA8/XA6/MN2/a_324_n18# AVSS 0.01fF
C625 XA20/XA1/MN5/a_324_n18# XA20/XA1/MN4/a_324_n18# 0.01fF
C626 XA3/XA11/MP1/S XA3/CEO 0.02fF
C627 AVDD XB1/XA3/MP0/a_216_334# 0.15fF
C628 XA0/XA4/A XA0/XA4/MP1/a_216_n18# 0.15fF
C629 XA2/CN0 EN 0.08fF
C630 XA7/EN XA6/XA1/XA1/MP0/a_216_n18# 0.01fF
C631 XA1/XA2/A XA1/XA1/XA5/MN2/S 0.05fF
C632 XA3/XA1/XA1/MP3/G XA3/XA1/XA1/MN2/S 0.08fF
C633 XA5/XA5/MN0/a_324_n18# XA5/XA4/A 0.07fF
C634 XA3/CN0 XA20/CNO 0.05fF
C635 XA7/XA1/XA5/MP1/S XA20/CNO 0.01fF
C636 XA5/XA5/MP1/a_216_n18# VREF 0.02fF
C637 XA4/XA1/XA5/MN1/S AVDD 0.02fF
C638 XA1/XA6/MP1/a_216_n18# XA1/CN0 0.15fF
C639 XA20/XA3a/MP0/a_216_n18# XA20/XA3a/MP1/a_216_n18# 0.01fF
C640 SARN CK_SAMPLE 0.02fF
C641 XA7/XA4/MN1/a_324_n18# XA7/XA4/MN2/a_324_n18# 0.01fF
C642 XA4/XA4/A XA4/XA4/MN3/a_324_n18# 0.15fF
C643 XA6/XA5/MP2/a_216_n18# XA6/CN0 0.01fF
C644 XA8/XA3/MP2/a_216_n18# VREF 0.03fF
C645 XA6/XA4/A AVSS 1.11fF
C646 XB1/XA3/MN0/a_324_n18# XB1/XA0/MN0/a_324_n18# 0.01fF
C647 XA5/XA6/MN1/S CK_SAMPLE 0.05fF
C648 XA5/XA1/XA4/MP2/S XA5/XA1/XA4/MP1/S 0.04fF
C649 XA0/CEIN XB1/XA4/MN1/S 0.01fF
C650 XB2/CKN SAR_IN 0.23fF
C651 XA1/XA4/MP1/a_216_n18# XA1/XA4/MP2/a_216_n18# 0.01fF
C652 XA3/CP0 XA3/XA4/MN1/a_324_n18# 0.03fF
C653 VREF D<8> 0.77fF
C654 XA2/XA6/MN1/S D<6> 0.01fF
C655 XA0/CEIN CK_SAMPLE_BSSW 4.95fF
C656 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC32a<0>/XRES8/B 0.02fF
C657 XB1/CKN XB1/XA4/MP1/a_216_n18# 0.08fF
C658 XA6/EN XA5/XA4/A 0.12fF
C659 XA8/EN XA7/XA1/XA4/MP1/S 0.02fF
C660 XA2/XA5/MP1/a_216_n18# VREF 0.02fF
C661 XA3/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C662 XA2/EN XA1/XA1/XA1/MP2/a_216_n18# 0.02fF
C663 XA1/XA11/A XA1/XA9/Y 0.14fF
C664 XA0/XA9/MP0/a_216_n18# AVDD 0.09fF
C665 XA4/XA1/XA4/MP0/a_216_n18# EN 0.07fF
C666 XB2/M6/a_324_n18# XA0/CEIN 0.15fF
C667 XA4/XA1/XA2/Y XA4/XA1/XA5/MN1/S 0.05fF
C668 XB1/M7/a_324_n18# XB1/M8/a_324_n18# 0.01fF
C669 XA2/XA4/A VREF 0.37fF
C670 XA0/CP1 XA2/CN1 0.12fF
C671 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128b<2>/XRES16/B 0.03fF
C672 XA6/XA11/MN0/a_324_n18# XA6/XA11/MN1/a_324_n18# 0.01fF
C673 XA2/XA5/MN2/a_324_n18# AVSS 0.01fF
C674 XA8/XA1/XA2/Y XA8/XA1/XA5/MN1/S 0.05fF
C675 XA3/XA11/MN1/a_324_n18# XA3/XA12/MN0/a_324_n18# 0.01fF
C676 XA5/XA1/XA1/MN0/a_324_n18# XA5/EN 0.09fF
C677 XA2/XA6/MN3/S AVSS 0.13fF
C678 XA8/XA1/XA5/MN2/a_324_n18# XA8/XA2/MN0/a_324_n18# 0.01fF
C679 XA4/XA2/MP0/a_216_n18# AVDD 0.08fF
C680 XA4/XA11/MP1/S VREF 0.01fF
C681 XA0/XA2/MP3/a_216_n18# XA0/XA2/MP2/a_216_n18# 0.01fF
C682 XA1/XA12/A XA1/XA9/B 0.01fF
C683 XA7/XA1/XA5/MP2/S XA7/XA4/A 0.02fF
C684 XA20/XA9/Y AVSS 1.58fF
C685 XA5/XA9/Y XA5/XA11/MN0/a_324_n18# 0.07fF
C686 XA2/XA1/XA1/MP2/S XA2/XA1/XA1/MP3/G 0.04fF
C687 XA1/CEO AVSS 0.64fF
C688 XA7/CP0 VREF 0.77fF
C689 XA4/XA1/XA4/MN1/S XA20/CPO 0.03fF
C690 CK_SAMPLE XA8/XA6/MN2/a_324_n18# 0.15fF
C691 XA6/XA4/MP0/a_216_n18# AVDD 0.08fF
C692 XB1/M4/G XB1/XA1/Y 0.12fF
C693 XA2/XA6/MN3/S XA2/XA9/B 0.09fF
C694 XA7/XA13/MN1/a_324_n18# AVSS 0.09fF
C695 XA5/XA9/MN0/a_324_n18# XA5/XA8/MN0/a_324_n18# 0.01fF
C696 XA8/XA1/XA2/Y XA8/XA1/XA4/MN0/a_324_n18# 0.02fF
C697 XA3/XA9/B AVDD 0.79fF
C698 XB1/M4/G XB1/CKN 0.28fF
C699 XDAC2/XC0/XRES1A/B SARN 1.51fF
C700 XA5/XA11/A XA5/XA11/MN0/a_324_n18# 0.09fF
C701 XDAC2/XC64b<1>/XRES8/B SARN 11.94fF
C702 XA8/XA4/MP2/a_216_n18# AVDD 0.07fF
C703 XA1/EN XA1/CN0 0.10fF
C704 VREF XA7/XA3/MP0/a_216_n18# 0.02fF
C705 XA4/CN1 VREF 0.76fF
C706 XDAC2/XC128b<2>/XRES1B/B AVSS 2.95fF
C707 XA1/CEO XA2/XA9/B 0.02fF
C708 XA0/XA1/XA4/MN1/a_324_n18# XA0/XA1/XA2/Y 0.09fF
C709 XA20/XA13/MN1/a_324_n18# XA20/XA13/MN1/a_324_334# 0.01fF
C710 XA6/XA1/XA4/MP2/S EN 0.03fF
C711 XA7/XA1/XA5/MN1/S XA20/CNO 0.02fF
C712 XA8/XA1/XA5/MP0/a_216_n18# XA8/XA1/XA5/MP1/a_216_n18# 0.01fF
C713 XA3/XA9/Y XA3/XA9/B 0.15fF
C714 XA20/XA2/MP1/a_216_n18# XA20/XA2/MP2/a_216_n18# 0.01fF
C715 D<3> XA5/XA1/XA1/MN2/S 0.01fF
C716 XA20/XA9/A XA20/XA12/Y 0.07fF
C717 XA20/XA9/A AVSS 2.26fF
C718 XA7/XA1/XA4/MN1/S XA7/XA1/XA4/MN2/S 0.04fF
C719 XA6/EN VREF 1.22fF
C720 XDAC2/XC128b<2>/XRES1B/B XDAC2/XC128a<1>/XRES1B/B 0.03fF
C721 XA5/XA4/MP2/a_216_n18# AVDD 0.07fF
C722 XA6/XA4/A EN 0.10fF
C723 XA20/XA3/MN1/a_324_n18# XA20/XA9/Y 0.07fF
C724 XA20/XA4/MP5_DMY/a_216_n18# XA20/XA4/MP6_DMY/a_216_n18# 0.01fF
C725 AVDD XB1/XA1/Y 0.45fF
C726 XA2/CN1 XA2/XA1/XA5/MN2/S 0.01fF
C727 XA6/XA12/A AVSS 0.42fF
C728 XA5/XA12/A VREF 0.03fF
C729 XA3/XA1/XA1/MP3/S XA20/CPO 0.01fF
C730 XA20/XA4/MP0/a_216_n18# XA20/XA4/MP0/a_216_334# 0.01fF
C731 XA0/CP1 D<7> 0.80fF
C732 XB1/XA5b/MN1/a_324_n18# AVSS 0.12fF
C733 AVDD XB1/CKN 1.81fF
C734 XA20/XA1/MP3_DMY/a_216_n18# AVDD 0.24fF
C735 XA2/XA6/MN2/a_324_n18# AVSS 0.01fF
C736 XB1/XCAPB1/XCAPB4/m3_252_308# XB1/XA4/GNG 0.13fF
C737 XA6/XA1/XA5/MP2/S XA6/XA2/A 0.06fF
C738 XB2/XA7/MP1/a_216_334# XB2/XA5/MP1/a_216_n18# 0.01fF
C739 XA4/XA2/MP2/a_216_n18# XA4/XA2/MP3/a_216_n18# 0.01fF
C740 XA4/XA6/MP3/S VREF 0.02fF
C741 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MN3/a_324_n18# 0.08fF
C742 AVDD XA1/CN1 1.39fF
C743 D<5> AVSS 3.42fF
C744 SAR_IN XA0/CEIN 0.34fF
C745 XA2/XA6/MN3/S CK_SAMPLE 0.03fF
C746 XA6/XA3/MN2/a_324_n18# XA6/XA4/A 0.01fF
C747 XDAC2/XC1/XRES4/B XDAC2/XC64a<0>/XRES8/B 0.01fF
C748 XA6/XA3/MN0/a_324_n18# XA6/XA2/A 0.07fF
C749 XA8/XA11/MP0/a_216_n18# XA8/XA11/A 0.07fF
C750 XA0/XA3/MP0/a_216_n18# D<8> 0.07fF
C751 XA2/XA3/MP2/a_216_n18# XA2/XA3/MP3/a_216_n18# 0.01fF
C752 XA5/XA13/MN1/a_324_334# XA5/XA13/MN1/a_324_n18# 0.01fF
C753 XA3/EN XA2/XA1/XA5/MP2/S 0.02fF
C754 XA7/XA9/B XA7/XA9/MN0/a_324_n18# 0.01fF
C755 XA20/XA2/MN2/a_324_n18# XA20/XA2/MN3/a_324_n18# 0.01fF
C756 XA20/XA9/Y CK_SAMPLE 0.03fF
C757 XA3/XA12/A XA2/CEO 0.18fF
C758 XA6/CN0 D<1> 0.05fF
C759 XA1/XA1/XA5/MN2/S XA1/CN1 0.01fF
C760 XA8/XA4/MP1/a_216_n18# XA8/XA4/A 0.15fF
C761 XDAC2/XC0/XRES2/B AVSS 3.67fF
C762 XA1/XA9/MP1/a_216_334# XA1/XA9/B 0.08fF
C763 XA20/CPO XA0/XA1/XA2/Y 0.21fF
C764 XA2/XA12/MN0/a_324_n18# XA2/XA11/MN1/a_324_n18# 0.01fF
C765 XA3/XA6/MP1/a_216_n18# AVDD 0.08fF
C766 XA8/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C767 XA4/XA1/XA5/MN2/S XA4/XA1/XA5/MP2/S 0.01fF
C768 XA3/XA1/XA1/MN2/S AVSS 0.27fF
C769 XA2/EN XA1/XA1/XA1/MP3/G 0.26fF
C770 XA2/XA1/XA1/MN1/a_324_n18# XA2/XA1/XA1/MN2/a_324_n18# 0.01fF
C771 XA20/XA9/Y EN 0.04fF
C772 XA5/XA9/MP1/a_216_n18# AVDD 0.09fF
C773 XA8/XA1/XA1/MP3/S XA8/XA1/XA1/MP3/G 0.04fF
C774 XA8/XA4/MP3/a_216_n18# VREF 0.02fF
C775 XA5/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C776 SARN XA20/XA4/MN5/a_324_n18# 0.15fF
C777 XA3/XA8/MP0/a_216_n18# XA3/XA9/A 0.07fF
C778 XA4/XA1/XA1/MP3/a_216_n18# AVDD 0.08fF
C779 XA6/XA9/Y XA6/XA12/A 0.02fF
C780 XA4/XA4/MN1/a_324_n18# XA4/XA4/MN0/a_324_n18# 0.01fF
C781 XA7/XA4/A XA8/XA2/A 0.03fF
C782 XA1/XA8/MP0/a_216_n18# AVDD 0.09fF
C783 XA3/XA4/MN0/a_324_n18# XA3/CN1 0.07fF
C784 XA4/XA13/MP1/a_216_n18# AVDD 0.13fF
C785 XA4/CP0 AVSS 0.91fF
C786 XA8/XA13/MN1/a_324_n18# AVSS 0.09fF
C787 XDAC1/XC64b<1>/XRES1A/B XDAC1/X16ab/XRES16/B 0.04fF
C788 XB1/XA3/MP0/S XB1/XA4/GNG 0.02fF
C789 XDAC1/XC32a<0>/XRES16/B XDAC1/XC128a<1>/XRES16/B 0.41fF
C790 XA2/CP0 XA2/XA5/MN1/a_324_n18# 0.15fF
C791 XA0/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C792 XA1/XA13/MN1/a_324_n18# XA1/XA12/A 0.07fF
C793 XA20/XA9/A CK_SAMPLE 0.10fF
C794 XA3/XA1/XA5/MN2/S AVSS 0.09fF
C795 XA7/CEO AVDD 0.77fF
C796 XB1/XA0/MN0/a_324_n18# AVSS 0.08fF
C797 AVDD XA0/XA1/XA1/MP0/a_216_n18# 0.15fF
C798 SARN SAR_IP 0.67fF
C799 XA5/CEO XA5/XA11/MP1/S 0.02fF
C800 XDAC2/X16ab/XRES1A/B XDAC2/X16ab/XRES8/B 0.12fF
C801 XDAC2/X16ab/XRES2/B XDAC2/X16ab/XRES4/B 0.55fF
C802 XDAC2/XC32a<0>/C1A AVSS 0.01fF
C803 XA1/CEO XA2/XA12/A 0.14fF
C804 XA4/XA1/XA1/MP3/a_216_n18# XA4/XA1/XA2/MP0/a_216_n18# 0.01fF
C805 XA5/XA3/MN3/a_324_n18# XA5/XA4/A 0.01fF
C806 XA3/CN1 XA3/XA4/A 0.61fF
C807 XA0/CP1 VREF 1.73fF
C808 XA2/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C809 XA20/XA11/Y VREF 0.01fF
C810 XA3/XA1/XA1/MP3/G AVDD 0.62fF
C811 XDAC1/XC128b<2>/XRES16/B XDAC1/XC128b<2>/XRES4/B 0.25fF
C812 XA4/XA13/MP1/a_216_n18# XA4/XA13/MP1/a_216_334# 0.01fF
C813 XA2/XA3/MP2/a_216_n18# D<6> 0.01fF
C814 XB1/M3/a_324_n18# XB1/M4/a_324_n18# 0.01fF
C815 XA6/CN0 XA3/CN1 0.05fF
C816 XDAC1/XC64b<1>/XRES1B/B AVSS 2.95fF
C817 XA0/XA12/MP0/a_216_n18# AVDD 0.08fF
C818 D<5> CK_SAMPLE 0.10fF
C819 XDAC1/XC128b<2>/XRES2/B SARP 3.05fF
C820 XA7/XA1/XA1/MP3/G XA7/XA1/XA1/MN3/a_324_n18# 0.08fF
C821 AVDD XA8/XA6/MP0/a_216_n18# 0.08fF
C822 XA7/CP0 XA8/CP0 0.03fF
C823 XA20/XA3/MN3/a_324_n18# SARN 0.15fF
C824 XA4/EN XA2/CN1 0.03fF
C825 XA8/XA6/MN0/a_324_n18# XA8/XA5/MN3/a_324_n18# 0.01fF
C826 XB2/M5/a_324_n18# XB2/M4/a_324_n18# 0.01fF
C827 XDAC1/XC32a<0>/XRES2/B XDAC1/XC128a<1>/XRES16/B 0.01fF
C828 D<4> XA0/CN0 0.07fF
C829 XA2/XA6/MP0/a_216_n18# VREF 0.01fF
C830 XDAC1/XC32a<0>/XRES1B/B AVSS 2.96fF
C831 XA1/DONE AVDD 0.21fF
C832 XDAC1/XC64b<1>/XRES1B/B XDAC1/X16ab/XRES1B/B 0.03fF
C833 D<5> EN 0.04fF
C834 XA6/CN0 D<2> 2.33fF
C835 XDAC1/XC64a<0>/XRES2/B XDAC1/XC64a<0>/XRES1A/B 0.25fF
C836 XA0/CP1 XA0/XA7/MP0/a_216_n18# 0.08fF
C837 XDAC1/XC64b<1>/XRES4/B XDAC1/XC64b<1>/XRES8/B 2.60fF
C838 XA7/XA2/MP2/a_216_n18# VREF 0.03fF
C839 XA1/XA1/XA1/MN2/S XA1/XA1/XA1/MP3/G 0.08fF
C840 XA20/XA9/MP0/a_216_334# AVDD 0.09fF
C841 XA1/XA1/XA5/MP2/S VREF 0.03fF
C842 XA3/XA3/MN3/a_324_n18# D<5> 0.02fF
C843 XA7/XA11/A XA7/CEO 0.05fF
C844 XA20/XA9/Y XA20/XA1/MN6/a_324_n18# 0.08fF
C845 AVDD XA20/XA3a/MP3/a_216_n18# 0.09fF
C846 AVDD XA8/XA9/MP1/a_216_n18# 0.09fF
C847 XA2/XA2/A XA3/EN 0.10fF
C848 XA6/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C849 XA6/CN0 XA7/CN0 3.63fF
C850 XA2/XA4/MP0/a_216_n18# AVDD 0.08fF
C851 XA5/CEO XA6/XA11/A 0.08fF
C852 XDAC1/XC128a<1>/XRES1B/B AVSS 2.95fF
C853 XA3/XA1/XA4/MP1/S EN 0.02fF
C854 XA2/CN0 XA2/CN1 1.69fF
C855 XA7/XA9/B AVDD 0.79fF
C856 XA4/CP0 CK_SAMPLE 0.09fF
C857 XA6/XA1/XA2/Y D<2> 0.02fF
C858 XA5/CEO XA6/CEO 0.04fF
C859 XA0/XA1/XA4/MN2/a_324_n18# XA0/XA1/XA2/Y 0.08fF
C860 XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MP3/S 0.04fF
C861 XA2/CP0 XA0/CN0 0.07fF
C862 XA4/XA4/MP0/a_216_n18# AVDD 0.08fF
C863 XA6/CN0 D<3> 0.13fF
C864 XA1/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C865 XA4/XA13/MN1/a_324_334# AVSS 0.10fF
C866 XB1/M5/a_324_n18# XB1/M4/a_324_n18# 0.01fF
C867 XA7/EN XA6/XA1/XA1/MN2/S 0.06fF
C868 XDAC1/XC32a<0>/XRES4/B XDAC1/XC32a<0>/XRES8/B 2.60fF
C869 XA2/XA4/A XA2/XA4/MP2/a_216_n18# 0.15fF
C870 XA2/XA6/MP3/a_216_n18# XA2/XA7/MP0/a_216_n18# 0.01fF
C871 XA20/XA4/MN2/a_324_n18# XA20/XA4/MN1/a_324_n18# 0.01fF
C872 XA20/XA11/MN1/a_324_n18# DONE 0.08fF
C873 XA4/XA13/MP1/a_216_n18# XA4/XA12/MP0/a_216_n18# 0.01fF
C874 XA4/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C875 EN XA2/XA1/XA5/MP0/a_216_n18# 0.16fF
C876 XA1/XA1/XA2/Y XA1/XA1/XA4/MN1/S 0.05fF
C877 XA0/XA9/A AVSS 0.29fF
C878 XA8/XA11/A XA8/XA9/Y 0.14fF
C879 XA6/XA6/MP2/a_216_n18# AVDD 0.09fF
C880 XA2/CN1 SARN 0.15fF
C881 XA6/XA4/MP3/a_216_n18# VREF 0.03fF
C882 XA3/XA1/XA5/MN2/S EN 0.02fF
C883 XDAC2/XC128b<2>/XRES16/B XA1/CN0 0.01fF
C884 AVDD XA2/XA11/A 0.45fF
C885 XA6/XA4/MN3/a_324_n18# XA6/XA5/MN0/a_324_n18# 0.01fF
C886 XB2/M4/G SARN 0.25fF
C887 XA7/XA1/XA1/MP3/S AVDD 0.13fF
C888 XA5/XA9/MN1/a_324_n18# XA5/XA9/B 0.09fF
C889 XA5/CN1 D<4> 0.01fF
C890 XA0/XA1/XA5/MN1/S XA0/XA1/XA2/Y 0.05fF
C891 XA3/XA2/MP2/a_216_n18# VREF 0.03fF
C892 XDAC2/XC128a<1>/XRES1A/B XDAC2/XC32a<0>/XRES8/B 0.03fF
C893 XA4/XA1/XA1/MP3/a_216_n18# XA5/EN 0.02fF
C894 XA1/XA13/MN1/a_324_n18# XA1/XA13/MN1/a_324_334# 0.01fF
C895 XA6/XA9/B XA6/XA6/MN1/S 0.05fF
C896 XA7/XA11/A XA7/XA9/B 0.02fF
C897 XDAC2/XC128a<1>/XRES16/B XA1/CN0 0.01fF
C898 XA5/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C899 XDAC2/XC0/XRES2/B XDAC2/XC0/XRES1A/B 0.25fF
C900 XA4/XA2/A XA4/CN1 0.57fF
C901 XA3/CP0 XA3/CN1 0.20fF
C902 XA8/XA1/XA4/MN1/S XA20/CNO 0.01fF
C903 XA6/XA1/XA5/MN2/S XA6/XA1/XA5/MP2/S 0.01fF
C904 XA8/XA12/A XA8/XA13/MP1/a_216_n18# 0.08fF
C905 XA4/XA1/XA4/MN1/S XA4/XA1/XA4/MP1/S 0.01fF
C906 XA7/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C907 XA8/XA4/MP3/a_216_n18# XA8/CP0 0.02fF
C908 XDAC1/XC64b<1>/XRES4/B XDAC1/XC0/XRES1A/B 0.01fF
C909 XDAC1/XC1/XRES16/B XDAC1/XC1/XRES4/B 0.25fF
C910 XA6/XA6/MP3/a_216_n18# XA6/XA6/MP2/a_216_n18# 0.01fF
C911 XA2/EN XA1/XA4/A 0.12fF
C912 XA1/XA8/MP0/a_216_n18# XA1/XA9/A 0.07fF
C913 XA6/EN XA4/XA2/A 0.03fF
C914 XA8/CEO XA20/XA12/MN0/a_324_n18# 0.08fF
C915 XB1/M4/G AVSS 0.96fF
C916 D<2> XA3/CP0 0.03fF
C917 XA0/CP0 XA0/XA2/A 0.03fF
C918 XA4/XA8/MP0/a_216_n18# XA4/XA9/MP0/a_216_n18# 0.01fF
C919 XA4/XA11/MP1/a_216_n18# XA4/XA11/A 0.08fF
C920 XA3/EN XA2/XA1/XA2/MN0/a_324_n18# 0.09fF
C921 XA20/CNO XA2/XA1/XA2/Y 0.22fF
C922 XA3/XA1/XA4/MN2/a_324_n18# XA3/EN 0.08fF
C923 XA8/CN0 XA8/XA5/MP2/a_216_n18# 0.01fF
C924 XA6/XA12/MP0/a_216_n18# XA6/XA12/A 0.07fF
C925 XA4/XA1/XA1/MN2/S XA4/EN 0.05fF
C926 XA7/CN0 XA3/CP0 0.04fF
C927 XA2/EN XA0/CP0 0.04fF
C928 XA2/XA2/MN1/a_324_n18# XA2/XA2/MN0/a_324_n18# 0.01fF
C929 XA20/XA2/N2 XA20/XA3/CO 0.03fF
C930 XA6/CN0 XA8/EN 0.04fF
C931 XDAC1/XC0/XRES16/B XA1/CN1 0.04fF
C932 XA3/XA5/MP3/a_216_n18# XA3/XA5/MP2/a_216_n18# 0.01fF
C933 XA1/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C934 XDAC2/XC64b<1>/XRES2/B AVSS 3.71fF
C935 XA0/XA2/A XA0/XA2/MN1/a_324_n18# 0.15fF
C936 XDAC2/XC32a<0>/XRES2/B AVSS 3.96fF
C937 XA20/XA3/MN1/a_324_n18# XA20/XA3/MN0/a_324_n18# 0.01fF
C938 D<6> D<4> 0.33fF
C939 XA8/XA1/XA5/MP2/S EN 0.03fF
C940 XA3/EN XA2/XA1/XA1/MP1/a_216_n18# 0.02fF
C941 XA5/XA1/XA1/MP3/S AVDD 0.13fF
C942 XDAC2/XC128b<2>/XRES8/B SARN 11.94fF
C943 XB2/XA3/B AVDD 2.43fF
C944 XA1/XA1/XA2/Y XA20/CPO 0.24fF
C945 XA3/XA5/MN2/a_324_n18# XA3/XA5/MN1/a_324_n18# 0.01fF
C946 XA6/XA1/XA4/MP1/a_216_n18# XA6/XA1/XA4/MP2/a_216_n18# 0.01fF
C947 XA0/XA9/A CK_SAMPLE 0.02fF
C948 XA4/XA2/MN0/a_324_n18# XA4/XA1/XA5/MN2/a_324_n18# 0.01fF
C949 XDAC2/XC128a<1>/XRES8/B XDAC2/XC32a<0>/XRES1B/B 0.02fF
C950 XB1/XA5/MP1/a_216_n18# XB1/XA4/GNG 0.01fF
C951 XA3/XA1/XA4/MN2/a_324_n18# XA3/XA1/XA4/MN1/a_324_n18# 0.01fF
C952 XA1/XA6/MN2/a_324_n18# AVSS 0.01fF
C953 D<3> XA3/CP0 0.01fF
C954 XA7/XA12/A VREF 0.03fF
C955 XA1/XA6/MP3/S AVDD 0.16fF
C956 XB2/M7/a_324_n18# XA0/CEIN 0.15fF
C957 D<7> SARN 0.03fF
C958 AVDD AVSS 42.85fF
C959 XA20/XA12/Y AVDD 0.86fF
C960 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128a<1>/XRES1A/B 0.03fF
C961 XA4/XA9/B XA3/CEO 0.02fF
C962 XA6/XA1/XA4/MN2/S XA6/EN 0.02fF
C963 XA5/XA3/MP3/a_216_n18# XA5/XA4/MP0/a_216_n18# 0.01fF
C964 XB2/XA5/MN1/a_324_n18# AVSS 0.09fF
C965 XB2/XA2/MP0/G XB2/XA5/MP1/a_216_n18# 0.08fF
C966 XA5/XA1/XA4/MN2/a_324_n18# XA5/XA1/XA2/Y 0.08fF
C967 XA1/XA3/MP0/a_216_n18# VREF 0.02fF
C968 XA20/XA1/MP4_DMY/a_216_n18# AVDD 0.24fF
C969 XA8/XA8/MN0/a_324_n18# XA8/XA9/A 0.09fF
C970 D<0> XA8/XA3/MN1/a_324_n18# 0.02fF
C971 XA1/XA9/A XA1/DONE 0.07fF
C972 XA6/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C973 XA20/XA3a/A XA20/XA3/CO 1.45fF
C974 XA4/XA2/MP3/a_216_n18# VREF 0.03fF
C975 XA5/XA4/MN2/a_324_n18# AVSS 0.01fF
C976 XA1/XA1/XA5/MN2/S AVSS 0.09fF
C977 XA4/EN VREF 1.19fF
C978 XA1/XA2/A XA1/CN1 0.62fF
C979 XA3/XA1/XA2/Y XA3/EN 0.14fF
C980 AVDD XA20/XA3a/MP2/a_216_n18# 0.08fF
C981 XA3/XA9/Y AVSS 0.22fF
C982 XA5/XA9/MP0/a_216_n18# AVDD 0.09fF
C983 XA6/XA9/Y XA6/XA9/MP1/a_216_334# 0.07fF
C984 XDAC1/XC128b<2>/XRES16/B AVSS 16.02fF
C985 XA2/CP0 D<6> 6.18fF
C986 XA20/XA11/MP0/a_216_n18# XA20/XA10/MP1/a_216_n18# 0.01fF
C987 XB1/CKN XB1/XA3/MP0/a_216_334# 0.09fF
C988 XA4/XA5/MP2/a_216_n18# VREF 0.03fF
C989 XA5/XA9/B AVDD 0.79fF
C990 XA20/XA3/MN5/a_324_n18# XA20/XA3/N1 0.01fF
C991 XA8/XA6/MN2/a_324_n18# XA8/XA6/MN3/a_324_n18# 0.01fF
C992 EN XA2/XA1/XA5/MP2/a_216_n18# 0.16fF
C993 XA2/XA9/B AVDD 0.79fF
C994 XB1/XA3/MP2/a_216_n18# XB1/XA3/B 0.02fF
C995 XA4/XA1/XA2/Y AVSS 0.30fF
C996 AVDD XA20/XA4/MP4_DMY/a_216_n18# 0.24fF
C997 XA6/CEO XA6/XA13/MP1/a_216_n18# 0.01fF
C998 XA8/EN XA7/XA8/MN0/a_324_n18# 0.06fF
C999 XA4/XA6/MP2/a_216_n18# XA4/XA6/MP3/a_216_n18# 0.01fF
C1000 XA4/XA6/MN3/S AVDD 0.01fF
C1001 XA1/CP0 XDAC1/XC128a<1>/XRES16/B 0.01fF
C1002 XA6/CN1 XA5/CN1 0.10fF
C1003 XA20/CPO XA0/XA1/XA1/MP3/G 0.14fF
C1004 D<4> SARP 0.06fF
C1005 XA4/XA1/XA2/Y XA4/XA1/XA5/MN1/a_324_n18# 0.09fF
C1006 SARN XA20/XA4/MN1/a_324_n18# 0.09fF
C1007 XA4/XA9/MN1/S AVSS 0.15fF
C1008 XA6/XA13/MN1/a_324_334# AVSS 0.10fF
C1009 XA3/XA1/XA4/MN1/a_324_n18# XA3/XA1/XA2/Y 0.09fF
C1010 XA2/CN0 VREF 0.69fF
C1011 XA6/XA9/Y AVDD 0.58fF
C1012 XA20/XA4/MN2/a_324_n18# XA20/XA4/MP0/S 0.01fF
C1013 XA1/XA9/MN1/S AVSS 0.15fF
C1014 XA0/XA4/MP0/a_216_n18# D<8> 0.08fF
C1015 XA3/XA1/XA4/MN0/a_324_n18# XA3/XA1/XA2/Y 0.02fF
C1016 XA7/XA11/A AVSS 0.27fF
C1017 XA0/XA1/XA1/MP3/a_216_n18# XA1/EN 0.02fF
C1018 XA8/XA1/XA4/MP2/S XA20/CPO 0.01fF
C1019 XA1/XA4/MN0/a_324_n18# XA1/XA4/MN1/a_324_n18# 0.01fF
C1020 XA20/XA9/Y XA20/XA2/MN0/a_324_n18# 0.14fF
C1021 XA7/XA1/XA4/MP1/S XA7/XA1/XA2/Y 0.01fF
C1022 XA20/XA4/MP6_DMY/a_216_n18# XA20/XA9/MP0/a_216_n18# 0.01fF
C1023 XA6/XA5/MP3/a_216_n18# XA6/CP0 0.15fF
C1024 EN XA2/XA1/XA4/MP0/a_216_n18# 0.07fF
C1025 XA4/XA3/MP2/a_216_n18# VREF 0.03fF
C1026 XA1/XA4/MP0/a_216_n18# XA1/XA3/MP3/a_216_n18# 0.01fF
C1027 XA2/XA2/MP1/a_216_n18# XA2/XA2/MP2/a_216_n18# 0.01fF
C1028 XDAC1/XC128b<2>/XRES4/B XDAC1/XC128b<2>/XRES1B/B 1.64fF
C1029 XA4/XA3/MP0/a_216_n18# XA4/XA3/MP1/a_216_n18# 0.01fF
C1030 XA8/XA3/MN2/a_324_n18# XA8/XA3/MN1/a_324_n18# 0.01fF
C1031 XA4/XA7/MN0/a_324_n18# XA5/EN 0.08fF
C1032 XA20/CPO D<8> 0.14fF
C1033 XA8/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C1034 XB1/XA3/B XB1/XA3/MN2/a_324_n18# 0.01fF
C1035 XA6/XA9/A XA5/XA9/A 0.02fF
C1036 XA1/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C1037 XDAC2/X16ab/XRES4/B XDAC2/X16ab/XRES16/B 0.25fF
C1038 XA3/XA2/MP2/a_216_n18# XA3/XA2/A 0.15fF
C1039 XA6/XA7/MP0/a_216_n18# XA7/EN 0.07fF
C1040 XA6/XA4/A XA5/XA4/A 0.16fF
C1041 XA2/CP0 SARP 0.07fF
C1042 XB2/XA1/MP0/G SARN 0.01fF
C1043 XDAC1/XC1/XRES1B/B XDAC1/XC64a<0>/XRES1A/B 0.63fF
C1044 XA20/XA2a/MN1/a_324_n18# XA20/XA3/CO 0.15fF
C1045 AVDD CK_SAMPLE 6.47fF
C1046 XA2/XA3/MN1/a_324_n18# XA2/XA3/MN2/a_324_n18# 0.01fF
C1047 XA8/XA2/MN2/a_324_n18# XA8/XA2/A 0.15fF
C1048 XA4/XA4/MP2/a_216_n18# XA4/XA4/MP1/a_216_n18# 0.01fF
C1049 XA7/CN0 XA7/XA5/MP2/a_216_n18# 0.01fF
C1050 XB2/M8/a_324_334# XA0/CEIN 0.09fF
C1051 XA4/XA6/MN1/S AVDD 0.01fF
C1052 XA2/XA4/A XA20/CPO 0.03fF
C1053 XA8/XA1/XA4/MP2/S XA8/XA1/XA4/MN2/S 0.01fF
C1054 XA7/XA2/MN2/a_324_n18# XA7/XA2/A 0.15fF
C1055 XA8/XA1/XA1/MN1/a_324_n18# XA8/XA1/XA1/MN2/a_324_n18# 0.01fF
C1056 XA8/XA2/MP3/a_216_n18# XA8/XA2/A 0.15fF
C1057 XA6/EN XA5/XA1/XA1/MP2/a_216_n18# 0.02fF
C1058 XB2/XA1/Y XB2/XA4/GNG 0.03fF
C1059 XA0/XA12/MN0/a_324_n18# XA0/XA13/MN1/a_324_n18# 0.01fF
C1060 XA4/XA3/MP1/a_216_n18# D<4> 0.03fF
C1061 XA20/CNO XA5/XA1/XA5/MN1/a_324_n18# 0.07fF
C1062 XA6/XA1/XA1/MP1/a_216_n18# AVDD 0.08fF
C1063 XA7/XA2/MP3/a_216_n18# AVDD 0.07fF
C1064 XA7/XA11/MN0/a_324_n18# XA7/XA11/A 0.09fF
C1065 XA2/XA9/MP1/a_216_n18# XA2/XA9/MP0/a_216_n18# 0.01fF
C1066 XB2/XA4/MN0/a_324_n18# XB2/XA4/MN1/a_324_n18# 0.01fF
C1067 XA6/XA1/XA5/MP0/a_216_n18# EN 0.16fF
C1068 XA1/CN0 XA0/CN0 6.53fF
C1069 XA2/XA1/XA1/MN2/a_324_n18# XA2/XA1/XA1/MN3/a_324_n18# 0.01fF
C1070 XA5/XA12/MP0/a_216_n18# XA5/XA11/MP1/a_216_n18# 0.01fF
C1071 XDAC2/XC128a<1>/XRES4/B XDAC2/XC128a<1>/XRES1A/B 0.29fF
C1072 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC64a<0>/XRES1A/B 0.01fF
C1073 XDAC1/XC1/XRES2/B AVSS 3.64fF
C1074 EN AVDD 25.90fF
C1075 XA3/XA4/MP2/a_216_n18# XA3/XA4/A 0.15fF
C1076 XA3/XA1/XA4/MN2/S XA3/EN 0.02fF
C1077 XA7/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C1078 XA2/XA5/MP3/a_216_n18# VREF 0.02fF
C1079 XA6/XA11/MN0/a_324_n18# XA6/XA9/MN1/a_324_334# 0.01fF
C1080 XA1/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C1081 XA20/XA2a/MP1/a_216_n18# XA20/XA2/MP6/a_216_334# 0.01fF
C1082 XA1/XA1/XA5/MN2/S EN 0.02fF
C1083 XA7/XA1/XA1/MN0/a_324_n18# XA7/XA1/XA1/MN1/a_324_n18# 0.01fF
C1084 XA8/XA1/XA1/MN2/S AVDD 0.07fF
C1085 D<5> XA2/CN1 0.05fF
C1086 XA6/XA11/MP0/a_216_n18# XA6/XA11/A 0.07fF
C1087 XB2/XA1/Y SAR_IN 0.04fF
C1088 XB2/XCAPB1/XCAPB0/m3_9756_132# XB2/XA4/GNG 0.02fF
C1089 XB1/XCAPB1/XCAPB0/m3_9828_132# XB1/XA3/B 0.21fF
C1090 AVDD XA8/XA6/MP3/a_216_n18# 0.08fF
C1091 XA20/XA4/MP4_DMY/a_216_n18# XA20/XA4/MP3_DMY/a_216_n18# 0.01fF
C1092 XA4/XA8/MN0/a_324_n18# XA5/EN 0.06fF
C1093 D<1> XA7/XA6/MN1/S 0.01fF
C1094 XA4/XA4/MP2/a_216_n18# VREF 0.03fF
C1095 XA8/XA12/MP0/a_216_n18# AVDD 0.08fF
C1096 XB1/XA1/MP0/G XB1/XA2/MP0/G 0.02fF
C1097 XA1/XA3/MP0/a_216_n18# XA1/XA2/MP3/a_216_n18# 0.01fF
C1098 XA0/XA1/XA2/MN0/a_324_n18# XA1/EN 0.09fF
C1099 XA6/XA1/XA4/MP1/S XA6/XA1/XA2/Y 0.01fF
C1100 XA4/XA1/XA2/Y EN 0.07fF
C1101 AVDD XA2/XA12/A 0.44fF
C1102 XA5/EN AVSS 1.25fF
C1103 XA0/XA4/A XA0/XA4/MN3/a_324_n18# 0.15fF
C1104 XB1/XA3/MP0/a_216_n18# XB1/XA3/B 0.01fF
C1105 AVDD XA8/XA6/MN3/S 0.01fF
C1106 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC64b<1>/XRES4/B 1.64fF
C1107 XDAC2/XC64b<1>/XRES2/B XDAC2/XC64b<1>/XRES8/B 1.58fF
C1108 XDAC1/XC128a<1>/XRES1B/B XDAC1/XC128b<2>/XRES8/B 0.02fF
C1109 XB1/CKN XB1/XA1/Y 0.08fF
C1110 XA3/XA1/XA1/MP3/S XA3/XA1/XA1/MP2/S 0.04fF
C1111 XDAC1/X16ab/XRES4/B XDAC1/X16ab/XRES16/B 0.25fF
C1112 XA1/XA11/MN1/a_324_n18# AVSS 0.01fF
C1113 XA2/XA2/MP1/a_216_n18# AVDD 0.08fF
C1114 XA1/XA9/A AVSS 0.31fF
C1115 XA1/XA1/XA2/Y XA1/CP0 0.01fF
C1116 XDAC2/XC128b<2>/XRES1B/B XDAC2/XC128b<2>/XRES8/B 0.12fF
C1117 XA2/XA7/MP0/a_216_n18# AVDD 0.09fF
C1118 XA6/XA1/XA5/MP1/S XA7/EN 0.02fF
C1119 XA1/XA4/MP1/a_216_n18# XA1/XA4/MP0/a_216_n18# 0.01fF
C1120 XA6/EN XA20/CPO 0.74fF
C1121 XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MP2/a_216_n18# 0.01fF
C1122 XA8/XA2/MP1/a_216_n18# XA8/XA2/A 0.15fF
C1123 XA3/XA2/A XA4/EN 0.10fF
C1124 XA7/XA4/MN2/a_324_n18# XA7/XA4/A 0.15fF
C1125 XA6/XA4/A VREF 0.37fF
C1126 XA0/CP1 XDAC1/XC64b<1>/XRES16/B 0.05fF
C1127 XA7/XA5/MN0/a_324_n18# XA7/XA5/MN1/a_324_n18# 0.01fF
C1128 XA4/XA9/A AVDD 0.62fF
C1129 XA8/XA4/A XA20/CNO 0.14fF
C1130 XA4/CP0 XA4/XA5/MP0/a_216_n18# 0.07fF
C1131 XA5/XA1/XA5/MN2/S XA20/CNO 0.01fF
C1132 XA8/CN1 AVDD 1.37fF
C1133 XA5/XA4/A XA5/XA4/MN1/a_324_n18# 0.15fF
C1134 XA8/XA12/A XA8/CEO 0.06fF
C1135 XA0/CP0 XDAC1/X16ab/XRES16/B 0.03fF
C1136 XA2/XA9/B XA1/XA9/A 0.02fF
C1137 XA7/XA5/MP0/a_216_n18# XA7/XA4/MP3/a_216_n18# 0.01fF
C1138 XA6/XA9/B XA6/XA6/MP1/S 0.07fF
C1139 XA20/XA2/MP5/a_216_n18# AVDD 0.10fF
C1140 XA6/XA11/MN1/a_324_n18# XA6/XA12/A 0.01fF
C1141 XA1/CN0 XA1/XA5/MP1/a_216_n18# 0.02fF
C1142 XDAC1/XC1/XRES4/B XDAC1/XC1/XRES1A/B 0.29fF
C1143 XA7/XA9/MN1/a_324_334# XA7/XA9/B 0.07fF
C1144 XA7/XA1/XA4/MP1/a_216_n18# XA7/XA1/XA4/MP2/a_216_n18# 0.01fF
C1145 XA7/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C1146 SARN XA20/XA4/MP0/S 0.19fF
C1147 XA2/CN1 XDAC2/XC32a<0>/C1A 0.04fF
C1148 XA7/XA11/MP1/a_216_n18# AVDD 0.08fF
C1149 XA5/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C1150 XA1/XA1/XA4/MN2/S XA1/EN 0.02fF
C1151 XDAC1/XC64a<0>/XRES1A/B SARP 1.50fF
C1152 XA2/CP0 XA2/XA4/MN1/a_324_n18# 0.03fF
C1153 XA4/XA1/XA4/MN1/a_324_n18# XA4/XA1/XA4/MN0/a_324_n18# 0.01fF
C1154 XA3/XA2/MP1/a_216_n18# XA3/CN1 0.02fF
C1155 D<3> XA5/XA3/MP3/a_216_n18# 0.02fF
C1156 XA4/XA9/B D<4> 0.05fF
C1157 XA6/CN1 XA7/EN 0.10fF
C1158 XDAC2/XC64b<1>/XRES4/B XDAC2/XC0/XRES16/B 0.03fF
C1159 XB2/XCAPB1/XCAPB0/m3_252_308# XB2/XA3/B 0.02fF
C1160 D<5> D<7> 0.79fF
C1161 XA7/XA2/A AVSS 0.28fF
C1162 XA4/XA9/Y XA4/XA12/A 0.02fF
C1163 XA20/XA9/Y VREF 0.07fF
C1164 XA4/EN XA3/XA1/XA2/MN0/a_324_n18# 0.09fF
C1165 XA4/CN0 D<4> 2.26fF
C1166 XA1/CEO VREF 0.05fF
C1167 XA5/EN CK_SAMPLE 0.09fF
C1168 XA20/XA3/N2 SARN 0.10fF
C1169 XA0/XA5/MN0/a_324_n18# XA0/XA4/MN3/a_324_n18# 0.01fF
C1170 XDAC1/XC0/XRES16/B AVSS 15.94fF
C1171 XA20/XA9/A XA20/XA4/MN1/a_324_n18# 0.07fF
C1172 D<6> XA1/CN0 0.04fF
C1173 XB2/XA3/B XB2/XA5b/MP1/a_216_n18# 0.02fF
C1174 XB2/M4/G XB2/M4/a_324_n18# 0.15fF
C1175 XA6/XA12/MP0/a_216_n18# AVDD 0.08fF
C1176 XA20/XA4/MN3/a_324_n18# XA20/XA4/MP0/S 0.01fF
C1177 XA6/EN XA5/XA1/XA4/MP0/a_216_n18# 0.08fF
C1178 XB1/XA4/MP0/a_216_n18# XB1/XA4/GNG 0.02fF
C1179 XB1/XCAPB1/XCAPB0/m3_324_308# XB1/XA3/B 0.02fF
C1180 AVDD XA8/XA9/MN1/S 0.01fF
C1181 XB1/CKN XB1/XA3/MN0/a_324_n18# 0.09fF
C1182 SAR_IP XB1/M4/G 0.62fF
C1183 XDAC2/XC32a<0>/XRES16/B AVSS 17.65fF
C1184 XA1/CP0 D<8> 0.03fF
C1185 XA1/XA9/A CK_SAMPLE 0.02fF
C1186 XA5/CN0 D<4> 0.01fF
C1187 XA4/XA2/A XA4/XA2/MP3/a_216_n18# 0.15fF
C1188 XB2/XA5b/MP1/a_216_n18# AVSS 0.02fF
C1189 XA0/CP1 XA0/XA4/MP0/a_216_n18# 0.01fF
C1190 XA6/XA5/MP2/a_216_n18# XA6/XA5/MP1/a_216_n18# 0.01fF
C1191 XA1/XA4/A XA1/XA5/MP0/a_216_n18# 0.08fF
C1192 XA4/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C1193 XA4/XA2/A XA4/EN 0.06fF
C1194 XA0/XA12/A XA0/XA13/MN1/a_324_n18# 0.07fF
C1195 XA4/XA1/XA1/MN0/a_324_n18# XA4/EN 0.08fF
C1196 SARN XA20/XA4/MN0/a_324_n18# 0.02fF
C1197 XDAC2/X16ab/XRES1B/B AVSS 2.95fF
C1198 XA5/EN EN 1.03fF
C1199 XA8/XA8/MN0/a_324_n18# XA8/XA9/MN0/a_324_n18# 0.01fF
C1200 XA2/XA1/XA1/MP1/a_216_n18# XA2/XA1/XA1/MP2/a_216_n18# 0.01fF
C1201 XA5/XA5/MN1/a_324_n18# XA5/CN0 0.02fF
C1202 VREF XA3/XA5/MP0/a_216_n18# 0.02fF
C1203 XA7/XA11/MP1/a_216_n18# XA7/XA11/A 0.08fF
C1204 SARN XDAC2/XC32a<0>/XRES4/B 6.32fF
C1205 XDAC1/XC128b<2>/XRES1B/B AVSS 2.95fF
C1206 XA1/XA11/A XA1/XA9/B 0.02fF
C1207 XA4/XA12/A XA4/XA11/MN1/a_324_n18# 0.01fF
C1208 XA0/CP1 XA20/CPO 0.05fF
C1209 XA6/XA1/XA1/MN1/a_324_n18# AVSS 0.01fF
C1210 XA2/XA4/MP3/a_216_n18# AVDD 0.07fF
C1211 XA3/XA4/MP2/a_216_n18# XA3/XA4/MP1/a_216_n18# 0.01fF
C1212 XA20/XA1/MN3/a_324_n18# SARP 0.15fF
C1213 XDAC1/XC128b<2>/XRES16/B XDAC1/X16ab/XRES1A/B 0.04fF
C1214 XA0/XA1/XA4/MP1/a_216_n18# XA0/XA1/XA4/MP0/a_216_n18# 0.01fF
C1215 XA7/XA3/MN0/a_324_n18# XA7/CN1 0.10fF
C1216 XA20/XA9/A VREF 0.03fF
C1217 XA8/XA4/MN0/a_324_n18# XA8/XA4/A 0.09fF
C1218 XA1/XA12/MP0/a_216_n18# XA1/XA11/MP1/a_216_n18# 0.01fF
C1219 XA6/XA1/XA5/MN1/S XA6/XA1/XA2/Y 0.05fF
C1220 XA6/XA1/XA5/MP0/a_216_n18# XA6/XA1/XA5/MP1/a_216_n18# 0.01fF
C1221 XA5/XA3/MP0/a_216_n18# AVDD 0.08fF
C1222 XA1/XA2/A AVSS 0.23fF
C1223 VREF XA8/XA5/MP3/a_216_n18# 0.02fF
C1224 XDAC2/XC64a<0>/XRES8/B SARN 11.94fF
C1225 AVDD SAR_IP 0.11fF
C1226 XDAC1/XC128b<2>/XRES1B/B XDAC1/X16ab/XRES1B/B 0.03fF
C1227 XA6/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C1228 EN XA0/XA1/XA5/MP2/a_216_n18# 0.16fF
C1229 XA4/XA2/MP2/a_216_n18# AVDD 0.07fF
C1230 XA7/XA12/MN0/a_324_n18# XA6/CEO 0.07fF
C1231 D<5> XA3/XA3/MP1/a_216_n18# 0.02fF
C1232 XA4/XA9/Y XA4/XA11/A 0.14fF
C1233 XA20/XA11/MP1/a_216_n18# DONE 0.07fF
C1234 XA8/XA1/XA5/MP0/a_216_n18# EN 0.15fF
C1235 XA6/XA12/A VREF 0.03fF
C1236 XA5/DONE AVDD 0.21fF
C1237 XA1/CN0 SARP 0.02fF
C1238 XA6/XA2/MN0/a_324_n18# XA6/XA2/A 0.08fF
C1239 XA6/XA1/XA1/MN2/a_324_n18# XA6/XA1/XA1/MN3/a_324_n18# 0.01fF
C1240 XA4/XA1/XA5/MN1/S AVSS 0.12fF
C1241 D<6> XA3/EN 0.42fF
C1242 XA5/XA13/MP1/a_216_n18# XA5/XA12/MP0/a_216_n18# 0.01fF
C1243 XDAC1/XC128b<2>/XRES16/B XDAC1/XC128b<2>/XRES8/B 1.42fF
C1244 XA3/XA1/XA1/MN3/a_324_n18# XA3/XA1/XA1/MP3/G 0.08fF
C1245 XA4/CP0 XA4/XA4/MP1/a_216_n18# 0.02fF
C1246 D<5> VREF 1.73fF
C1247 XA1/XA4/A XA1/XA4/MP3/a_216_n18# 0.15fF
C1248 XA8/XA1/XA5/MN2/S XA8/XA4/A 0.02fF
C1249 XA4/XA12/MN0/a_324_n18# XA4/XA11/MN1/a_324_n18# 0.01fF
C1250 XDAC2/XC1/XRES1B/B XDAC2/XC64a<0>/XRES8/B 0.02fF
C1251 XA5/XA4/MP1/a_216_n18# XA5/XA4/MP0/a_216_n18# 0.01fF
C1252 XA4/XA1/XA1/MN1/a_324_n18# AVSS 0.01fF
C1253 XA3/XA1/XA4/MP2/a_216_n18# XA3/XA1/XA5/MP0/a_216_n18# 0.01fF
C1254 XA3/XA1/XA4/MP0/a_216_n18# XA3/XA1/XA2/MP0/a_216_n18# 0.01fF
C1255 XA5/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C1256 D<0> XA20/XA3/CO 0.01fF
C1257 XA7/XA2/MP3/a_216_n18# XA7/XA2/A 0.15fF
C1258 XA4/XA5/MP1/a_216_n18# XA4/XA5/MP0/a_216_n18# 0.01fF
C1259 XA8/XA1/XA1/MP2/a_216_n18# XA20/CPO 0.07fF
C1260 XDAC1/XC128a<1>/XRES8/B AVSS 9.08fF
C1261 XB2/XA3/MN2/a_324_n18# XB2/XA3/MN1/a_324_n18# 0.01fF
C1262 XA4/XA9/A XA5/EN 0.09fF
C1263 AVDD XA6/XA1/XA1/MP3/G 0.63fF
C1264 XA2/XA13/MP1/a_216_n18# XA2/XA12/MP0/a_216_n18# 0.01fF
C1265 XA8/XA4/MN1/a_324_n18# XA8/CP0 0.03fF
C1266 EN XA7/XA2/A 0.11fF
C1267 XA1/CN0 XA1/XA5/MP3/a_216_n18# 0.02fF
C1268 XA8/XA1/XA4/MN1/S XA8/XA4/A 0.02fF
C1269 XA8/XA9/MN1/a_324_334# XA8/XA9/Y 0.09fF
C1270 XA4/XA11/A XA4/XA11/MN1/a_324_n18# 0.07fF
C1271 XA0/XA2/A XA0/XA1/XA2/Y 0.01fF
C1272 XA1/XA1/XA4/MN2/S XA1/XA1/XA4/MP2/S 0.01fF
C1273 XB2/CKN XB2/XA4/MP0/a_216_n18# 0.15fF
C1274 XA8/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C1275 XB2/XA3/B XDAC2/XC1/XRES1A/B 0.21fF
C1276 D<3> XA5/XA1/XA2/Y 0.02fF
C1277 XA2/XA1/XA1/MP3/a_216_n18# XA2/XA1/XA2/MP0/a_216_n18# 0.01fF
C1278 XB2/XA3/MN0/a_324_n18# XB2/XA3/MN1/a_324_n18# 0.01fF
C1279 XA0/XA6/MP1/S XA0/CN0 0.02fF
C1280 XB2/XA7/MN1/a_324_334# XB2/XA5/MN1/a_324_n18# 0.01fF
C1281 D<6> XA2/XA1/XA1/MN2/S 0.02fF
C1282 XA20/XA9/Y XA20/XA4/MP0/S 0.05fF
C1283 XA4/EN XA3/XA1/XA1/MP3/a_216_n18# 0.01fF
C1284 XA20/XA11/MN0/a_324_n18# XA20/XA11/MN1/a_324_n18# 0.01fF
C1285 XDAC2/XC1/XRES1A/B AVSS 2.78fF
C1286 XDAC1/XC0/XRES2/B XDAC1/XC0/XRES16/B 1.61fF
C1287 XDAC1/XC1/XRES16/B XDAC1/XC64a<0>/XRES16/B 0.41fF
C1288 XA4/CP0 VREF 0.77fF
C1289 XB2/M4/G XB1/M4/G 0.07fF
C1290 XA0/XA1/XA4/MN1/S XA20/CPO 0.03fF
C1291 XA5/XA5/MP0/a_216_n18# AVDD 0.08fF
C1292 XA7/XA1/XA4/MP1/a_216_n18# XA7/XA1/XA4/MP0/a_216_n18# 0.01fF
C1293 XB1/XA3/MN1/a_324_n18# XB1/XA3/MN2/a_324_n18# 0.01fF
C1294 XA2/XA1/XA2/Y XA2/XA1/XA5/MN2/a_324_n18# 0.07fF
C1295 XA7/XA9/MN1/a_324_334# XA7/XA11/MN0/a_324_n18# 0.01fF
C1296 XA7/XA1/XA5/MP1/S XA7/XA1/XA5/MP2/S 0.04fF
C1297 XA3/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C1298 XA5/XA3/MP3/a_216_n18# XA5/XA3/MP2/a_216_n18# 0.01fF
C1299 XA2/CP0 XA2/XA5/MP2/a_216_n18# 0.15fF
C1300 XDAC1/XC64b<1>/XRES8/B XDAC1/XC64b<1>/XRES1A/B 0.12fF
C1301 XA7/CEO XA7/XA9/B 0.03fF
C1302 XA20/XA9/Y XA20/XA3/N2 0.03fF
C1303 XDAC2/XC64a<0>/XRES16/B XDAC2/XC64a<0>/XRES4/B 0.25fF
C1304 XA2/DONE XA2/XA9/Y 0.06fF
C1305 XDAC1/XC64b<1>/XRES4/B SARP 6.32fF
C1306 D<1> XA7/XA6/MP1/S 0.02fF
C1307 XA1/XA2/A EN 0.11fF
C1308 XA2/CN1 AVDD 1.41fF
C1309 XA3/XA9/B AVSS 0.61fF
C1310 XA0/XA1/XA5/MN1/S XA0/XA1/XA5/MN2/S 0.04fF
C1311 XA5/XA12/MP0/a_216_n18# XA4/CEO 0.08fF
C1312 XA8/XA2/MP0/a_216_n18# AVDD 0.08fF
C1313 XA4/XA5/MP0/a_216_n18# AVDD 0.08fF
C1314 XA0/XA13/MP1/a_216_n18# AVDD 0.13fF
C1315 XA6/XA6/MP0/a_216_n18# VREF 0.01fF
C1316 XA6/XA1/XA5/MN2/a_324_n18# XA6/EN 0.08fF
C1317 XA0/XA5/MN3/a_324_n18# XA0/XA6/MN0/a_324_n18# 0.01fF
C1318 XA20/XA9/A XA20/XA4/MP0/S 0.13fF
C1319 XA3/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C1320 XA20/XA9/Y XA8/CP0 0.02fF
C1321 XB2/M4/G AVDD 0.65fF
C1322 XDAC1/XC128a<1>/XRES16/B XDAC1/XC128a<1>/XRES2/B 1.61fF
C1323 XB2/CKN XB2/XA3/MP0/a_216_n18# 0.08fF
C1324 XA4/XA1/XA5/MP1/S XA4/XA4/A 0.02fF
C1325 XDAC2/XC0/XRES16/B XA0/CN0 0.02fF
C1326 XDAC1/XC32a<0>/XRES4/B SARP 6.32fF
C1327 XA1/XA3/MP1/a_216_n18# XA1/XA3/MP0/a_216_n18# 0.01fF
C1328 XA4/XA4/A XA3/XA4/A 0.16fF
C1329 XA2/XA1/XA1/MP3/G XA2/XA1/XA1/MP3/a_216_n18# 0.07fF
C1330 XA3/XA2/MP0/a_216_n18# AVDD 0.08fF
C1331 XB1/XCAPB1/XCAPB4/m3_9756_132# XB1/XA4/GNG 0.02fF
C1332 XA4/XA1/XA5/MN1/S EN 0.01fF
C1333 XA5/XA1/XA4/MN2/S XA20/CNO 0.01fF
C1334 XDAC2/XC64b<1>/XRES16/B XDAC2/X16ab/XRES8/B 0.03fF
C1335 XA20/XA13/MN1/a_324_334# AVDD 0.01fF
C1336 XA8/XA3/MN0/a_324_n18# XA8/CN1 0.10fF
C1337 XA20/XA3a/MN1/a_324_n18# XA20/XA3a/MN0/a_324_n18# 0.01fF
C1338 XB1/XA1/Y AVSS 0.33fF
C1339 XA20/XA9/Y XA20/XA9/MN0/a_324_n18# 0.08fF
C1340 XA20/XA3/MP3/a_216_n18# XA20/XA3a/A 0.01fF
C1341 XA20/XA9/A XA20/XA3/N2 0.07fF
C1342 XA20/CNO XA2/XA1/XA4/MN2/S 0.01fF
C1343 XA3/XA1/XA5/MN0/a_324_n18# XA3/EN 0.07fF
C1344 XDAC1/XC128a<1>/XRES4/B SARP 6.32fF
C1345 XA20/CNO XA3/XA1/XA1/MP2/a_216_n18# 0.08fF
C1346 XA5/XA1/XA1/MP3/G AVDD 0.62fF
C1347 XDAC2/XC64b<1>/XRES8/B XDAC2/X16ab/XRES1B/B 0.02fF
C1348 XB1/CKN AVSS 0.75fF
C1349 XDAC2/XC1/XRES16/B XDAC2/XC1/XRES2/B 1.61fF
C1350 XA0/CP0 XA3/CP0 0.61fF
C1351 XA2/XA8/MN0/a_324_n18# XA2/XA9/B 0.01fF
C1352 XA2/XA9/MP1/a_216_n18# XA2/XA9/MP1/a_216_334# 0.01fF
C1353 XA8/XA1/XA5/MP2/S VREF 0.03fF
C1354 SARP XB1/M3/a_324_n18# 0.01fF
C1355 XA6/CN0 XA6/XA2/A 0.04fF
C1356 XA2/XA4/A XA2/XA1/XA5/MP1/S 0.02fF
C1357 XA1/CN1 AVSS 2.61fF
C1358 XB1/XCAPB1/XCAPB2/m3_9828_132# XB1/XA3/B 0.21fF
C1359 XA6/XA1/XA4/MN2/S XA6/XA1/XA4/MP2/S 0.01fF
C1360 XA20/XA1/MP3_DMY/a_216_n18# XA20/XA1/MP4_DMY/a_216_n18# 0.01fF
C1361 XA0/CP1 XA1/CP0 0.10fF
C1362 XA2/XA9/B XA2/XA9/MN1/a_324_334# 0.07fF
C1363 SAR_IP XB1/M6/a_324_n18# 0.01fF
C1364 XDAC2/XC64b<1>/XRES1A/B XDAC2/X16ab/XRES1A/B 0.03fF
C1365 XA20/XA9/A XA20/XA4/MN0/a_324_n18# 0.08fF
C1366 XA0/XA4/MN2/a_324_n18# XA0/XA4/MN1/a_324_n18# 0.01fF
C1367 XA8/XA5/MP3/a_216_n18# XA8/CP0 0.15fF
C1368 D<1> XA7/XA3/MN3/a_324_n18# 0.02fF
C1369 XB1/XCAPB1/XCAPB2/m3_252_308# XB1/XA4/GNG 0.13fF
C1370 XA4/XA6/MP1/a_216_n18# XA4/CN0 0.15fF
C1371 XB1/XA3/MN2/a_324_n18# XB1/XA4/MN0/a_324_n18# 0.01fF
C1372 XA20/CNO XA6/XA1/XA1/MN2/S 0.03fF
C1373 XA5/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C1374 XA7/XA5/MP2/a_216_n18# XA7/XA5/MP1/a_216_n18# 0.01fF
C1375 XA7/XA2/MN3/a_324_n18# XA7/CN1 0.03fF
C1376 XA6/CN1 XA6/CP0 0.03fF
C1377 XA6/XA1/XA4/MN2/S XA6/XA4/A 0.06fF
C1378 XA1/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C1379 XA6/XA1/XA1/MP3/G XA6/XA1/XA1/MP3/a_216_n18# 0.07fF
C1380 D<5> XA3/XA2/A 0.06fF
C1381 XA6/XA2/A XA6/XA1/XA2/Y 0.01fF
C1382 XA1/CP0 XA1/XA4/MN3/a_324_n18# 0.02fF
C1383 XA0/XA9/A VREF 0.04fF
C1384 XA4/EN XA20/CPO 0.73fF
C1385 XA3/XA1/XA2/Y XA3/CN1 0.04fF
C1386 XDAC1/XC64b<1>/XRES1A/B XDAC1/XC0/XRES1A/B 0.03fF
C1387 XA6/XA9/A XA6/DONE 0.07fF
C1388 XB2/M8/a_324_n18# XA0/CEIN 0.15fF
C1389 D<1> XA7/XA4/A 0.26fF
C1390 VREF XA2/XA2/MP2/a_216_n18# 0.03fF
C1391 D<5> XA3/XA6/MN1/S 0.01fF
C1392 XDAC2/X16ab/XRES16/B XA1/CN0 0.01fF
C1393 XA4/XA2/MP0/a_216_n18# EN 0.08fF
C1394 XA5/XA4/A AVDD 1.42fF
C1395 XA20/XA9/A XA20/XA9/MN0/a_324_n18# 0.09fF
C1396 XA0/XA6/MP3/S XA1/EN 0.02fF
C1397 XA3/CN0 D<4> 0.06fF
C1398 XA3/XA9/B CK_SAMPLE 0.10fF
C1399 XA8/ENO XA20/XA3/CO 0.34fF
C1400 D<7> AVDD 1.85fF
C1401 AVDD XA8/XA9/B 0.79fF
C1402 XA7/XA5/MN1/a_324_n18# XA7/CP0 0.15fF
C1403 XA5/XA4/A XA5/XA4/MN2/a_324_n18# 0.15fF
C1404 XA1/CP0 XA1/XA5/MN3/a_324_n18# 0.15fF
C1405 XA4/CN0 XA1/CN0 0.10fF
C1406 XA5/XA1/XA4/MN2/a_324_n18# XA5/XA1/XA4/MN1/a_324_n18# 0.01fF
C1407 D<5> XA3/XA4/MP0/a_216_n18# 0.01fF
C1408 XA8/XA1/XA1/MP2/S AVDD 0.11fF
C1409 XA7/XA9/MP1/a_216_n18# AVDD 0.09fF
C1410 XA4/XA6/MP2/a_216_n18# AVDD 0.09fF
C1411 XA3/XA3/MP3/a_216_n18# VREF 0.03fF
C1412 XA4/XA5/MP1/a_216_n18# VREF 0.02fF
C1413 XA5/XA9/MP0/a_216_n18# XA5/XA9/MP1/a_216_n18# 0.01fF
C1414 SARP XB1/XA3/B 0.41fF
C1415 XA4/CN0 XA4/XA1/XA1/MP3/G 0.02fF
C1416 XA2/CN0 XA20/CPO 0.05fF
C1417 XA7/CN0 XA7/XA6/MP1/S 0.02fF
C1418 SARP XB1/M5/a_324_n18# 0.02fF
C1419 AVDD XA8/XA6/MP3/S 0.15fF
C1420 XA7/CEO AVSS 0.56fF
C1421 XDAC1/XC128b<2>/XRES4/B AVSS 5.49fF
C1422 XA5/XA9/MP1/a_216_n18# XA5/XA9/B 0.07fF
C1423 XB2/CKN SARN 0.04fF
C1424 XA5/CN0 XA1/CN0 0.11fF
C1425 XB1/XA3/MN0/a_324_n18# AVSS 0.01fF
C1426 XA1/XA1/XA1/MP3/G XA1/EN 0.09fF
C1427 XA1/XA6/MN1/a_324_n18# XA1/XA6/MN0/a_324_n18# 0.01fF
C1428 XA1/XA3/MN1/a_324_n18# XA1/CN1 0.16fF
C1429 XA5/XA5/MP2/a_216_n18# AVDD 0.07fF
C1430 XA3/XA9/B XA3/XA7/MN0/a_324_n18# 0.01fF
C1431 XA6/XA4/MN2/a_324_n18# XA6/XA4/A 0.15fF
C1432 XA5/XA2/MP1/a_216_n18# XA5/XA2/MP0/a_216_n18# 0.01fF
C1433 AVDD XA20/XA2a/MP2/a_216_n18# 0.08fF
C1434 XA4/XA4/MP1/a_216_n18# AVDD 0.07fF
C1435 XA0/XA5/MP1/a_216_n18# VREF 0.02fF
C1436 XDAC1/XC128b<2>/XRES1B/B XDAC1/X16ab/XRES1A/B 0.63fF
C1437 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128b<2>/XRES2/B 0.25fF
C1438 XA1/XA9/B XA1/XA6/MP1/S 0.07fF
C1439 XA3/CN0 XA2/CP0 0.03fF
C1440 XA4/XA1/XA1/MN2/S AVDD 0.05fF
C1441 XA2/XA9/Y XA2/XA11/MP0/a_216_n18# 0.08fF
C1442 XA6/XA9/A XA6/XA9/MP0/a_216_n18# 0.14fF
C1443 XA1/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C1444 XA3/XA1/XA1/MP3/G AVSS 0.11fF
C1445 XA3/XA2/A XA3/XA1/XA5/MN2/S 0.05fF
C1446 XA7/XA12/A XA7/XA9/Y 0.02fF
C1447 XA8/XA1/XA1/MP0/a_216_n18# XA8/XA1/XA1/MP1/a_216_n18# 0.01fF
C1448 XA20/CPO SARN 0.09fF
C1449 XA5/CN1 XA5/XA4/MP0/a_216_n18# 0.08fF
C1450 XA3/CN0 XA3/XA5/MP2/a_216_n18# 0.01fF
C1451 D<1> XA0/CN0 0.06fF
C1452 D<1> XA7/XA6/MP2/a_216_n18# 0.07fF
C1453 XDAC2/X16ab/XRES8/B SARN 11.94fF
C1454 XA4/XA2/A XA4/XA2/MN3/a_324_n18# 0.15fF
C1455 XA8/XA1/XA1/MP3/G XA20/CNO 0.06fF
C1456 XA20/CPO XA2/XA1/XA4/MN1/S 0.03fF
C1457 XA2/XA4/A XA2/XA1/XA5/MN1/S 0.02fF
C1458 XA5/EN XA5/XA1/XA5/MN0/a_324_n18# 0.07fF
C1459 XDAC1/XC128b<2>/XRES8/B XDAC1/XC128b<2>/XRES1B/B 0.12fF
C1460 XA3/XA3/MP1/a_216_n18# AVDD 0.07fF
C1461 XDAC1/XC64b<1>/XRES2/B XDAC1/X16ab/XRES2/B 0.05fF
C1462 XA1/DONE AVSS 0.15fF
C1463 EN XA1/CN1 0.07fF
C1464 XB2/XA5b/MN1/a_324_n18# AVDD 0.01fF
C1465 XA6/XA2/MP2/a_216_n18# VREF 0.03fF
C1466 XA1/XA7/MN0/a_324_n18# AVSS 0.01fF
C1467 XA4/XA9/B XA4/XA9/MN0/a_324_n18# 0.01fF
C1468 XDAC1/XC64b<1>/XRES8/B XDAC1/XC64b<1>/XRES2/B 1.58fF
C1469 XA5/CP0 D<4> 0.01fF
C1470 XA2/XA1/XA2/Y XA2/XA1/XA4/MN1/a_324_n18# 0.09fF
C1471 XA20/XA3/N1 SARN 0.33fF
C1472 XA4/XA2/MP1/a_216_n18# XA4/CN1 0.01fF
C1473 XA2/XA2/A XA2/XA2/MN3/a_324_n18# 0.15fF
C1474 VREF AVDD 68.61fF
C1475 XB2/XA1/MP0/G AVDD 0.28fF
C1476 D<2> XA7/XA4/A 0.01fF
C1477 XA5/CP0 XA5/XA5/MN1/a_324_n18# 0.15fF
C1478 XA7/XA2/MN2/a_324_n18# AVSS 0.01fF
C1479 XA2/EN XA1/XA1/XA2/Y 0.14fF
C1480 XA2/EN XA1/XA1/XA5/MP1/S 0.02fF
C1481 XA4/XA9/A XA3/XA9/B 0.02fF
C1482 XA6/XA1/XA4/MP1/S XA6/XA1/XA4/MN1/S 0.01fF
C1483 XDAC1/XC128a<1>/XRES1B/B XDAC1/XC128b<2>/XRES1A/B 0.63fF
C1484 XA7/XA9/B AVSS 0.61fF
C1485 VREF XA0/XA2/MP1/a_216_n18# 0.02fF
C1486 XA0/XA9/B XA0/XA9/MN0/a_324_n18# 0.01fF
C1487 XA5/XA5/MN3/a_324_n18# XA5/XA6/MN0/a_324_n18# 0.01fF
C1488 XA5/XA1/XA1/MP3/G XA5/EN 0.09fF
C1489 XA7/CN0 XA7/XA4/A 0.12fF
C1490 XA6/XA9/A XA6/XA11/A 0.01fF
C1491 XA20/XA3a/MP3/a_216_n18# XA20/XA3a/MP2/a_216_n18# 0.01fF
C1492 XA3/XA9/Y VREF 0.03fF
C1493 XA8/XA3/MP1/a_216_n18# D<0> 0.03fF
C1494 XB2/XCAPB1/XCAPB1/m3_9756_132# XB2/XA3/B 0.07fF
C1495 XA0/XA1/XA1/MN3/a_324_n18# XA0/XA1/XA1/MP3/G 0.08fF
C1496 XB2/XA7/MP1/a_216_334# AVDD 0.15fF
C1497 XA4/XA1/XA5/MP2/S XA4/XA4/A 0.02fF
C1498 XA6/XA12/MN0/a_324_n18# XA6/XA13/MN1/a_324_n18# 0.01fF
C1499 XA6/CN0 XA6/XA6/MP1/S 0.02fF
C1500 XA1/XA1/XA5/MN0/a_324_n18# XA1/EN 0.07fF
C1501 XA7/XA1/XA1/MP2/S AVDD 0.09fF
C1502 XA0/XA4/A XA0/XA4/MN0/a_324_n18# 0.09fF
C1503 XDAC2/XC0/XRES16/B SARP 0.03fF
C1504 XA8/XA11/MN0/a_324_n18# AVSS 0.01fF
C1505 XA0/XA7/MP0/a_216_n18# AVDD 0.09fF
C1506 XA2/XA1/XA2/Y XA2/XA1/XA4/MN2/S 0.05fF
C1507 XA3/XA13/MN1/a_324_n18# XA3/XA12/A 0.07fF
C1508 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128b<2>/XRES8/B 0.21fF
C1509 XA3/CN0 XA3/XA6/MP1/S 0.02fF
C1510 XA5/XA1/XA1/MP3/G XA5/XA1/XA2/MP0/a_216_n18# 0.08fF
C1511 XA3/CN1 XA0/CN0 0.39fF
C1512 EN XA0/XA1/XA1/MP0/a_216_n18# 0.06fF
C1513 XA4/XA7/MN0/a_324_n18# XA4/XA8/MN0/a_324_n18# 0.01fF
C1514 XA1/XA4/MN2/a_324_n18# AVSS 0.01fF
C1515 XA2/XA11/A AVSS 0.28fF
C1516 XA4/XA4/MN0/a_324_n18# XA4/XA3/MN3/a_324_n18# 0.01fF
C1517 XA7/XA1/XA1/MP3/S AVSS 0.02fF
C1518 XA1/XA1/XA4/MN2/a_324_n18# XA1/EN 0.08fF
C1519 XA5/XA4/A XA5/EN 0.20fF
C1520 XA7/XA11/A VREF 0.02fF
C1521 D<3> XA5/XA2/A 0.07fF
C1522 D<0> XA8/XA4/MP0/a_216_n18# 0.01fF
C1523 XA4/XA7/MN0/a_324_n18# AVSS 0.01fF
C1524 XA2/EN XA0/XA1/XA1/MP3/G 0.01fF
C1525 XA6/XA4/A XA20/CPO 0.03fF
C1526 XA20/CNO XA0/XA1/XA5/MN1/a_324_n18# 0.07fF
C1527 XA20/XA13/MP1/a_216_334# AVDD 0.17fF
C1528 XB2/XA3/MN1/a_324_n18# XB2/XA3/MP0/S 0.01fF
C1529 XA6/XA6/MP3/S D<2> 0.02fF
C1530 XA6/XA4/MN2/a_324_n18# XA6/XA4/MN1/a_324_n18# 0.01fF
C1531 XB2/XA7/MP1/a_216_n18# XB2/XA4/GNG 0.02fF
C1532 XA8/ENO XA8/XA1/XA2/MP0/a_216_n18# 0.08fF
C1533 XA8/XA1/XA2/Y AVDD 0.35fF
C1534 XA0/CP0 XDAC1/XC64a<0>/XRES16/B 0.05fF
C1535 XA3/XA8/MP0/a_216_n18# XA3/XA7/MP0/a_216_n18# 0.01fF
C1536 SARN XA0/CEIN 0.62fF
C1537 EN XA3/XA1/XA1/MP3/G 0.10fF
C1538 XA8/XA2/MN1/a_324_n18# XA8/XA2/MN2/a_324_n18# 0.01fF
C1539 D<2> XA0/CN0 0.09fF
C1540 XA3/XA5/MN2/a_324_n18# XA3/CP0 0.15fF
C1541 XA2/CN1 XDAC2/XC32a<0>/XRES16/B 0.04fF
C1542 XA8/CEO XA20/XA11/MP1/S 0.01fF
C1543 XA8/XA11/MP1/a_216_n18# XA8/XA11/MP0/a_216_n18# 0.01fF
C1544 XA7/XA11/MN1/a_324_n18# XA7/XA12/MN0/a_324_n18# 0.01fF
C1545 D<7> XA1/XA9/A 0.01fF
C1546 XA3/XA1/XA5/MN1/a_324_n18# XA3/XA1/XA5/MN2/a_324_n18# 0.01fF
C1547 XA0/CP1 XA0/XA6/MN1/S 0.01fF
C1548 XA1/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C1549 XA7/CEO XA8/XA12/MP0/a_216_n18# 0.08fF
C1550 XB1/XCAPB1/XCAPB3/m3_9828_132# XB1/XA4/GNG 0.04fF
C1551 XA0/XA2/A D<8> 0.62fF
C1552 XA20/XA9/MP0/a_216_334# CK_SAMPLE 0.01fF
C1553 XA2/XA9/B XA2/XA11/A 0.03fF
C1554 XA7/CN0 XA0/CN0 0.72fF
C1555 XA7/XA6/MP2/a_216_n18# XA7/CN0 0.08fF
C1556 XB2/XA4/GNG XB2/XCAPB1/XCAPB1/m3_9828_132# 0.04fF
C1557 XA2/XA6/MP1/a_216_n18# D<6> 0.01fF
C1558 XA4/XA3/MN2/a_324_n18# XA4/XA3/MN3/a_324_n18# 0.01fF
C1559 XA2/EN D<8> 0.03fF
C1560 XA1/CP0 XA1/XA5/MN1/a_324_n18# 0.15fF
C1561 XA2/XA3/MP0/a_216_n18# XA2/CN1 0.07fF
C1562 XA5/XA2/MP3/a_216_n18# XA5/XA2/A 0.15fF
C1563 XA1/XA9/B XA1/XA9/Y 0.15fF
C1564 XA2/XA4/A XA2/XA4/MN2/a_324_n18# 0.15fF
C1565 XA7/XA9/B CK_SAMPLE 0.10fF
C1566 XA4/XA2/A XA4/XA2/MN1/a_324_n18# 0.15fF
C1567 XA4/XA1/XA1/MN2/S XA5/EN 0.06fF
C1568 D<4> XA20/CNO 0.06fF
C1569 XA1/XA2/A XA2/CN1 0.04fF
C1570 D<3> XA0/CN0 0.14fF
C1571 XA5/XA12/A XA5/XA13/MN1/a_324_n18# 0.07fF
C1572 D<1> D<6> 0.04fF
C1573 XA2/EN XA2/XA4/A 0.14fF
C1574 XA8/XA3/MP0/a_216_n18# XA8/XA2/A 0.08fF
C1575 XA3/XA3/MP3/a_216_n18# XA3/XA4/MP0/a_216_n18# 0.01fF
C1576 XA20/XA9/Y XA20/CPO 0.10fF
C1577 XA6/XA8/MN0/a_324_n18# XA6/XA9/MN0/a_324_n18# 0.01fF
C1578 XA2/XA1/XA4/MN2/a_324_n18# XA2/XA1/XA5/MN0/a_324_n18# 0.01fF
C1579 XA8/XA2/A XA20/CNO 0.06fF
C1580 XA6/XA13/MP1/a_216_334# XA6/XA13/MP1/a_216_n18# 0.01fF
C1581 XA20/XA2/N2 SARP 0.04fF
C1582 XA5/XA1/XA5/MP2/S XA5/XA1/XA5/MN2/S 0.01fF
C1583 AVDD XA20/XA4/MP0/S 0.59fF
C1584 XA1/XA1/XA1/MN2/a_324_n18# XA1/XA1/XA1/MN1/a_324_n18# 0.01fF
C1585 XA1/XA4/A XA1/EN 0.20fF
C1586 XA5/XA1/XA1/MP3/S AVSS 0.02fF
C1587 XA5/XA11/A XA5/XA11/MP1/a_216_n18# 0.08fF
C1588 XB2/XA3/B AVSS 5.05fF
C1589 XA8/EN XA7/XA4/A 0.12fF
C1590 XA6/XA1/XA1/MP2/S AVDD 0.11fF
C1591 XA0/XA3/MP0/a_216_n18# AVDD 0.08fF
C1592 XA1/XA1/XA1/MP0/a_216_n18# XA1/XA1/XA1/MP1/a_216_n18# 0.01fF
C1593 XA20/XA3a/A XA20/XA2a/MP3/a_216_n18# 0.01fF
C1594 XA7/XA11/MP1/S XA6/CEO 0.02fF
C1595 XA2/EN XA1/XA8/MN0/a_324_n18# 0.06fF
C1596 XA0/XA9/MN1/a_324_n18# XA0/XA9/A 0.07fF
C1597 XA6/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C1598 XA1/XA2/MP3/a_216_n18# AVDD 0.07fF
C1599 XA20/XA12/Y AVSS 0.23fF
C1600 XA20/XA9/Y XA20/XA3/N1 0.22fF
C1601 XA20/XA3/MP4/a_216_n18# XA20/XA3a/A 0.07fF
C1602 XA0/CP0 XA1/EN 0.12fF
C1603 SAR_IP XB1/XA1/Y 0.04fF
C1604 XA2/CP0 XA20/CNO 0.05fF
C1605 XA1/CP0 SARN 0.03fF
C1606 XA4/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C1607 XA5/EN VREF 1.22fF
C1608 XA5/XA2/MN3/a_324_n18# XA5/XA2/A 0.15fF
C1609 XA1/XA5/MP2/a_216_n18# XA1/XA5/MP1/a_216_n18# 0.01fF
C1610 XA4/XA13/MN1/a_324_334# XA4/XA13/MN1/a_324_n18# 0.01fF
C1611 XA20/XA3/N2 AVDD 0.45fF
C1612 D<7> XDAC1/XC0/XRES16/B 0.01fF
C1613 XDAC2/XC128a<1>/XRES1B/B AVSS 2.95fF
C1614 SAR_IP XB1/CKN 0.21fF
C1615 XA5/XA1/XA5/MP1/a_216_n18# XA5/XA1/XA5/MP0/a_216_n18# 0.01fF
C1616 XDAC1/X16ab/XRES1B/B AVSS 2.95fF
C1617 XDAC2/XC128b<2>/XRES4/B XDAC2/X16ab/XRES4/B 0.10fF
C1618 XDAC2/XC128b<2>/XRES1B/B XDAC2/X16ab/XRES8/B 0.02fF
C1619 XA3/XA2/A AVDD 1.07fF
C1620 XA6/XA5/MP0/a_216_n18# VREF 0.02fF
C1621 XA3/DONE XA3/XA9/A 0.07fF
C1622 XA8/XA2/MN2/a_324_n18# XA8/XA2/MN3/a_324_n18# 0.01fF
C1623 XDAC1/XC128b<2>/XRES16/B XDAC1/XC128b<2>/XRES1A/B 1.60fF
C1624 XDAC2/XC32a<0>/XRES2/B XDAC2/XC32a<0>/XRES4/B 0.55fF
C1625 XA3/XA13/MP1/a_216_n18# XA3/XA13/MP1/a_216_334# 0.01fF
C1626 XA1/XA9/A VREF 0.04fF
C1627 XA6/XA4/MN3/a_324_n18# XA6/CP0 0.02fF
C1628 XA20/XA9/A XA20/CPO 0.14fF
C1629 XA3/XA6/MN1/S AVDD 0.01fF
C1630 XA20/XA2/MN2/a_324_n18# SARP 0.15fF
C1631 XA5/XA9/B AVSS 0.61fF
C1632 XDAC2/XC128a<1>/XRES16/B XDAC2/XC32a<0>/XRES8/B 0.03fF
C1633 XA6/XA1/XA5/MP1/S XA20/CNO 0.01fF
C1634 XA2/XA9/B AVSS 0.61fF
C1635 AVDD XA8/CP0 1.42fF
C1636 XA0/XA1/XA5/MN2/a_324_n18# XA0/XA1/XA5/MN1/a_324_n18# 0.01fF
C1637 XDAC2/XC0/XRES1B/B SARP 0.05fF
C1638 XA3/CN0 XA1/CN0 2.28fF
C1639 XDAC2/XC128a<1>/XRES2/B XDAC2/XC128a<1>/XRES4/B 0.55fF
C1640 D<1> SARP 0.09fF
C1641 XA4/XA6/MN3/S AVSS 0.13fF
C1642 XDAC1/X16ab/XRES2/B XDAC1/X16ab/XRES4/B 0.55fF
C1643 XA0/XA2/A XA0/XA2/MP0/a_216_n18# 0.08fF
C1644 XA5/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C1645 XDAC1/XC64b<1>/XRES8/B XDAC1/X16ab/XRES4/B 0.01fF
C1646 XA3/XA4/MP0/a_216_n18# AVDD 0.08fF
C1647 XA1/XA8/MN0/a_324_n18# XA1/XA9/MN0/a_324_n18# 0.01fF
C1648 XA5/CP0 XA5/XA5/MN2/a_324_n18# 0.15fF
C1649 XA1/XA1/XA1/MP3/a_216_n18# AVDD 0.08fF
C1650 D<6> XA3/CN1 0.13fF
C1651 D<3> XA5/CN1 0.43fF
C1652 XA6/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C1653 XA6/XA9/Y AVSS 0.22fF
C1654 XDAC1/XC128b<2>/XRES4/B XDAC1/X16ab/XRES1A/B 0.01fF
C1655 XA20/XA9/A XA20/XA3/N1 0.21fF
C1656 D<7> XA1/XA2/A 0.06fF
C1657 D<5> XA20/CPO 0.06fF
C1658 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC64b<1>/XRES16/B 0.12fF
C1659 XA2/XA12/A XA2/XA11/A 0.07fF
C1660 XA3/XA1/XA1/MP1/a_216_n18# AVDD 0.07fF
C1661 AVDD XA8/XA9/A 0.64fF
C1662 XA20/XA3/N1 XA20/XA2/MN4/a_324_n18# 0.01fF
C1663 AVDD XA20/XA4/MP5_DMY/a_216_n18# 0.24fF
C1664 XA2/XA3/MP1/a_216_n18# XA2/XA3/MP2/a_216_n18# 0.01fF
C1665 XA1/XA11/MN1/a_324_n18# XA1/XA11/MN0/a_324_n18# 0.01fF
C1666 D<2> D<6> 0.42fF
C1667 XA6/XA1/XA2/MP0/a_216_n18# XA6/XA1/XA4/MP0/a_216_n18# 0.01fF
C1668 XA3/XA1/XA4/MP1/S XA20/CPO 0.03fF
C1669 XA0/XA6/MP2/a_216_n18# XA0/CN0 0.08fF
C1670 XA20/XA1/MP6_DMY/a_216_n18# XA20/XA1/MP5_DMY/a_216_n18# 0.01fF
C1671 XA1/XA4/A XA2/XA2/A 0.03fF
C1672 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128b<2>/XRES16/B 1.60fF
C1673 XDAC1/XC128b<2>/XRES8/B XDAC1/XC128b<2>/XRES4/B 2.60fF
C1674 XA5/XA2/MP3/a_216_n18# XA5/CN1 0.02fF
C1675 CK_SAMPLE AVSS 4.54fF
C1676 XA20/XA12/Y CK_SAMPLE 0.17fF
C1677 XA1/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C1678 VREF XA7/XA2/A 0.36fF
C1679 XA5/XA2/A XA5/XA2/MP0/a_216_n18# 0.08fF
C1680 XA4/XA6/MN1/S AVSS 0.15fF
C1681 XA5/XA9/Y XA5/XA9/MN1/a_324_334# 0.09fF
C1682 XA1/XA4/A XA1/XA4/MP2/a_216_n18# 0.15fF
C1683 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC32a<0>/XRES16/B 0.12fF
C1684 XA2/XA4/A XA2/XA3/MN2/a_324_n18# 0.01fF
C1685 XA8/XA6/MN0/a_324_n18# XA8/XA6/MN1/a_324_n18# 0.01fF
C1686 D<1> XA7/EN 0.07fF
C1687 XA5/XA2/MP2/a_216_n18# XA5/XA2/MP1/a_216_n18# 0.01fF
C1688 XA1/XA9/B XA1/XA9/MP1/a_216_n18# 0.07fF
C1689 XA7/XA1/XA4/MN1/a_324_n18# XA7/XA1/XA2/Y 0.09fF
C1690 XA3/CN0 XA3/EN 0.10fF
C1691 XA7/XA9/MN0/a_324_n18# XA7/XA9/MN1/a_324_n18# 0.01fF
C1692 XA4/XA2/A AVDD 1.07fF
C1693 XA0/XA2/A XA0/XA1/XA5/MN2/S 0.05fF
C1694 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128a<1>/XRES16/B 0.04fF
C1695 XDAC2/XC64a<0>/XRES16/B XA1/CN0 0.16fF
C1696 XA2/XA1/XA5/MN2/S XA2/XA1/XA5/MN1/S 0.04fF
C1697 D<3> D<6> 0.04fF
C1698 XA1/XA4/A XA1/XA1/XA4/MP2/S 0.05fF
C1699 XA8/XA1/XA5/MN2/S XA8/XA2/A 0.05fF
C1700 EN AVSS 2.87fF
C1701 XB2/XA4/GNG XB2/XCAPB1/XCAPB3/m3_252_308# 0.13fF
C1702 XA3/CN1 SARP 0.05fF
C1703 XA7/XA1/XA5/MN2/S AVDD 0.02fF
C1704 SARP XB1/XA1/MP0/G 0.01fF
C1705 XDAC1/XC0/XRES2/B AVSS 3.67fF
C1706 XB2/XA0/MN0/a_324_n18# AVSS 0.08fF
C1707 XA2/XA4/MP2/a_216_n18# AVDD 0.07fF
C1708 XA5/XA9/B CK_SAMPLE 0.08fF
C1709 XA2/XA9/B CK_SAMPLE 0.09fF
C1710 XA4/XA7/MN0/a_324_n18# XA4/XA6/MN3/a_324_n18# 0.01fF
C1711 XA20/XA9/A XA20/XA9/MP0/a_216_n18# 0.07fF
C1712 XA1/XA1/XA5/MP1/a_216_n18# XA1/XA1/XA5/MP2/a_216_n18# 0.01fF
C1713 XA3/XA4/MN2/a_324_n18# XA3/XA4/MN1/a_324_n18# 0.01fF
C1714 XA8/XA5/MN0/a_324_n18# XA8/CP0 0.09fF
C1715 XA3/XA7/MN0/a_324_n18# AVSS 0.01fF
C1716 XA0/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C1717 XA4/XA6/MN3/S CK_SAMPLE 0.03fF
C1718 XA8/XA12/A XA8/XA11/A 0.07fF
C1719 XA20/XA1/MN5/a_324_n18# SARP 0.16fF
C1720 XA20/XA2/MN1/a_324_n18# XA20/XA2/MN2/a_324_n18# 0.01fF
C1721 XA20/XA1/MN1/a_324_n18# XA20/XA1/MN2/a_324_n18# 0.01fF
C1722 XDAC2/XC0/XRES8/B SARN 12.03fF
C1723 XA2/CN1 XA1/CN1 4.91fF
C1724 XB1/XA1/MP0/G XB1/XA4/MN1/a_324_334# 0.08fF
C1725 XA8/XA1/XA1/MN2/S AVSS 0.30fF
C1726 XA2/XA3/MP0/a_216_n18# VREF 0.02fF
C1727 XA6/XA3/MN2/a_324_n18# AVSS 0.01fF
C1728 XA5/CP0 XA5/XA4/MP3/a_216_n18# 0.02fF
C1729 D<2> SARP 0.05fF
C1730 XA4/XA2/A XA4/XA1/XA2/Y 0.01fF
C1731 XA7/XA1/XA4/MN1/S AVDD 0.02fF
C1732 XA3/XA6/MP0/a_216_n18# XA3/CP0 0.08fF
C1733 XA5/XA2/MN3/a_324_n18# XA5/CN1 0.03fF
C1734 XA0/CP1 XA0/XA2/A 0.05fF
C1735 XDAC1/XC64b<1>/XRES4/B XDAC1/XC0/XRES4/B 0.10fF
C1736 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC0/XRES8/B 0.02fF
C1737 XA1/XA2/A VREF 0.36fF
C1738 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC32a<0>/XRES2/B 0.23fF
C1739 XA2/XA12/A AVSS 0.42fF
C1740 XA7/CN0 SARP 0.02fF
C1741 XA7/XA12/MP0/a_216_n18# XA7/XA13/MP1/a_216_n18# 0.01fF
C1742 XA1/XA1/XA1/MP3/S AVDD 0.13fF
C1743 XA1/XA5/MP2/a_216_n18# XA1/XA5/MP3/a_216_n18# 0.01fF
C1744 XA6/XA1/XA4/MN2/S AVDD 0.02fF
C1745 AVSS XA8/XA6/MN3/S 0.12fF
C1746 XA2/EN XA0/CP1 0.02fF
C1747 D<1> XA7/XA3/MP1/a_216_n18# 0.03fF
C1748 XA0/XA1/XA1/MP3/S AVDD 0.14fF
C1749 XB2/XCAPB1/XCAPB4/m3_9828_132# XB2/XA3/B 0.21fF
C1750 XA1/XA6/MN3/a_324_n18# XA1/XA6/MN2/a_324_n18# 0.01fF
C1751 XA8/XA1/XA4/MP1/S XA8/XA1/XA4/MN1/S 0.01fF
C1752 XA6/XA1/XA5/MP2/S XA6/XA4/A 0.02fF
C1753 XA20/XA3/N2 XA20/XA3/MP2/a_216_n18# 0.01fF
C1754 XB2/XA2/MP0/G AVDD 0.45fF
C1755 XA4/XA3/MN0/a_324_n18# XA4/CN1 0.10fF
C1756 XA7/XA5/MP3/a_216_n18# XA7/XA6/MP0/a_216_n18# 0.01fF
C1757 XA20/XA10/MN1/a_324_n18# XA20/XA9/MN0/a_324_334# 0.01fF
C1758 XA0/XA9/Y XA0/XA9/A 0.04fF
C1759 XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MN3/a_324_n18# 0.08fF
C1760 XA2/CP0 XA2/XA5/MP0/a_216_n18# 0.07fF
C1761 D<3> SARP 0.07fF
C1762 XB2/XA2/MP0/G XB2/XA5/MN1/a_324_n18# 0.06fF
C1763 XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MP2/S 0.04fF
C1764 XB1/M2/a_324_n18# XB1/M1/a_324_n18# 0.01fF
C1765 XA4/XA9/A XA4/XA8/MN0/a_324_n18# 0.09fF
C1766 XDAC2/XC0/XRES1A/B AVSS 2.94fF
C1767 XA6/XA7/MN0/a_324_n18# AVSS 0.01fF
C1768 XDAC2/XC64b<1>/XRES8/B AVSS 9.08fF
C1769 XB1/XA5/MN1/a_324_n18# AVSS 0.09fF
C1770 XA2/XA9/B XA2/XA12/A 0.01fF
C1771 XA4/XA6/MN1/S CK_SAMPLE 0.05fF
C1772 AVDD XA2/XA1/XA1/MP0/a_216_n18# 0.15fF
C1773 XDAC1/XC64a<0>/XRES4/B XDAC1/XC64a<0>/XRES1A/B 0.29fF
C1774 XA1/CEO XA2/CEO 0.04fF
C1775 XA5/XA3/MN1/a_324_n18# XA5/XA3/MN0/a_324_n18# 0.01fF
C1776 XA2/CP0 XA2/XA1/XA2/Y 0.02fF
C1777 XA4/XA9/A AVSS 0.31fF
C1778 XA8/CN1 AVSS 0.82fF
C1779 XA0/XA4/MN2/a_324_n18# AVSS 0.01fF
C1780 XDAC2/XC128b<2>/XRES16/B XDAC2/XC128a<1>/XRES4/B 0.03fF
C1781 XA6/XA5/MP2/a_216_n18# XA6/CP0 0.15fF
C1782 XA5/XA4/MP2/a_216_n18# XA5/XA4/A 0.15fF
C1783 XA4/EN XA3/XA1/XA1/MP2/S 0.14fF
C1784 XA1/XA1/XA5/MP2/S XA2/EN 0.02fF
C1785 XA7/XA3/MN3/a_324_n18# XA7/CN1 0.15fF
C1786 D<2> XA7/EN 0.43fF
C1787 XA3/XA1/XA1/MP3/a_216_n18# AVDD 0.08fF
C1788 XA1/XA6/MP1/S XA1/CN0 0.02fF
C1789 AVDD XB1/XA7/MP1/a_216_334# 0.15fF
C1790 XA5/CN1 XA5/XA3/MP2/a_216_n18# 0.15fF
C1791 XA3/XA11/A XA3/CEO 0.04fF
C1792 XDAC1/XC1/XRES16/B XDAC1/XC1/XRES1B/B 0.12fF
C1793 XA7/XA4/MP0/a_216_n18# XA7/XA3/MP3/a_216_n18# 0.01fF
C1794 XB1/M4/G XB1/XA4/MN1/a_324_n18# 0.01fF
C1795 XA20/XA2/MP3/a_216_n18# XA20/XA2/MP4/a_216_n18# 0.01fF
C1796 XA1/XA3/MP2/a_216_n18# AVDD 0.07fF
C1797 XA7/CN0 XA7/EN 0.17fF
C1798 XDAC1/XC64b<1>/XRES1A/B SARP 1.50fF
C1799 XA6/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C1800 XDAC2/XC128a<1>/XRES4/B XDAC2/XC128a<1>/XRES16/B 0.25fF
C1801 XA3/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C1802 XA7/CN1 XA7/XA4/A 0.58fF
C1803 XB2/CKN XB2/XA4/MN0/a_324_n18# 0.09fF
C1804 D<7> XA1/CN1 0.89fF
C1805 XB1/XCAPB1/XCAPB3/m3_324_308# XB1/XA3/B 0.02fF
C1806 XA20/CNO XA1/CN0 0.05fF
C1807 XA0/XA12/MP0/a_216_n18# XA0/XA13/MP1/a_216_n18# 0.01fF
C1808 D<1> XA4/CN0 0.04fF
C1809 XA1/XA1/XA4/MN1/S AVDD 0.02fF
C1810 XA4/XA2/MN2/a_324_n18# XA4/CN1 0.02fF
C1811 XA6/EN XA5/XA1/XA1/MN2/S 0.12fF
C1812 XA4/CP0 XA4/XA4/MN3/a_324_n18# 0.02fF
C1813 XDAC1/XC0/XRES1A/B XDAC1/XC0/XRES1B/B 0.01fF
C1814 XA0/CP0 XA0/XA5/MP2/a_216_n18# 0.15fF
C1815 XA4/XA1/XA1/MP3/G XA20/CNO 0.06fF
C1816 XA20/XA10/MN1/S XA20/XA11/Y 0.07fF
C1817 D<5> XA1/CP0 0.24fF
C1818 CK_SAMPLE XA8/XA6/MN3/S 0.03fF
C1819 XA6/XA4/MP0/a_216_n18# VREF 0.02fF
C1820 AVSS XA8/XA9/MN1/S 0.15fF
C1821 XA5/XA9/Y XA4/CEO 0.03fF
C1822 XA5/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C1823 D<1> XA5/CN0 0.04fF
C1824 XA5/XA7/MP0/a_216_n18# XA5/XA8/MP0/a_216_n18# 0.01fF
C1825 XA4/XA2/A XA5/EN 0.10fF
C1826 XA7/XA5/MP0/a_216_n18# XA7/XA4/A 0.08fF
C1827 XDAC1/X16ab/XRES1A/B AVSS 2.95fF
C1828 XA7/XA1/XA1/MN2/S XA7/EN 0.05fF
C1829 XA6/XA1/XA0/MN1/a_324_n18# XA6/XA1/XA1/MN0/a_324_n18# 0.01fF
C1830 XA20/CPO XA2/XA1/XA4/MN0/a_324_n18# 0.09fF
C1831 XA3/XA9/B VREF 0.12fF
C1832 XA2/EN XA2/XA1/XA5/MN0/a_324_n18# 0.07fF
C1833 XA2/XA4/MP0/a_216_n18# XA2/CN1 0.08fF
C1834 XA8/XA4/MP2/a_216_n18# VREF 0.03fF
C1835 XA6/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C1836 XA1/XA3/MP1/a_216_n18# AVDD 0.07fF
C1837 XA6/XA2/MN0/a_324_n18# XA6/EN 0.07fF
C1838 XA0/XA9/Y AVDD 0.58fF
C1839 XB2/XA4/GNG XB2/XCAPB1/XCAPB2/m3_9828_132# 0.04fF
C1840 XDAC1/XC128b<2>/XRES1B/B XDAC1/XC128b<2>/XRES1A/B 0.01fF
C1841 XA20/XA3/N1 XA20/XA3/MN0/a_324_n18# 0.01fF
C1842 XA1/XA11/MN1/a_324_n18# XA1/XA12/MN0/a_324_n18# 0.01fF
C1843 XA0/XA9/B XA0/XA6/MP1/S 0.07fF
C1844 XA4/XA9/A CK_SAMPLE 0.02fF
C1845 XA6/XA2/MP3/a_216_n18# XA6/XA2/MP2/a_216_n18# 0.01fF
C1846 XDAC1/X16ab/XRES1A/B XDAC1/X16ab/XRES1B/B 0.01fF
C1847 XA5/XA11/A XA4/CEO 0.09fF
C1848 XA1/XA9/B XA2/XA9/A 0.02fF
C1849 XA6/XA1/XA4/MN1/a_324_n18# XA6/XA1/XA2/Y 0.09fF
C1850 XA1/XA2/A XA1/XA2/MP3/a_216_n18# 0.15fF
C1851 XA1/XA1/XA1/MP3/G XA1/XA1/XA1/MN3/a_324_n18# 0.08fF
C1852 XB1/XA3/B XB1/XA4/GNG 434.15fF
C1853 XA5/XA6/MN3/a_324_n18# XA5/XA6/MN2/a_324_n18# 0.01fF
C1854 XDAC2/XC64a<0>/XRES1B/B SARN 1.79fF
C1855 XDAC1/XC128b<2>/XRES8/B AVSS 9.08fF
C1856 XA4/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C1857 XA7/CEO XA8/XA9/B 0.02fF
C1858 XA6/XA2/MP3/a_216_n18# AVDD 0.07fF
C1859 XDAC2/X16ab/XRES16/B XA3/CN1 0.07fF
C1860 XA5/XA4/MP2/a_216_n18# VREF 0.03fF
C1861 SAR_IP AVSS 0.72fF
C1862 XB2/CKN AVDD 1.73fF
C1863 XA20/CNO XA3/EN 0.93fF
C1864 XA8/XA1/XA1/MN1/a_324_n18# XA20/CNO 0.07fF
C1865 XDAC2/XC32a<0>/XRES4/B XDAC2/XC32a<0>/XRES16/B 0.25fF
C1866 XA0/XA4/MP0/a_216_n18# AVDD 0.08fF
C1867 XA5/DONE AVSS 0.15fF
C1868 XA8/CN1 EN 0.02fF
C1869 XA4/CN0 XA3/CN1 0.15fF
C1870 VREF XA1/CN1 0.77fF
C1871 XA8/XA1/XA1/MP3/G XA8/XA1/XA2/MN0/a_324_n18# 0.06fF
C1872 XA6/CN0 D<8> 0.05fF
C1873 XDAC2/XC1/XRES1B/B XDAC2/XC64a<0>/XRES1B/B 0.03fF
C1874 XDAC2/XC64a<0>/XRES8/B XDAC2/XC32a<0>/XRES16/B 0.03fF
C1875 XA7/XA4/MP3/a_216_n18# XA7/CP0 0.02fF
C1876 XA20/CPO AVDD 8.27fF
C1877 XA8/EN XA7/EN 1.77fF
C1878 XA2/XA4/A XA3/XA4/A 0.03fF
C1879 XA5/CN0 XA3/CN1 0.05fF
C1880 XA6/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C1881 XB2/XA1/Y SARN 0.02fF
C1882 XA3/XA9/A XA4/EN 0.09fF
C1883 D<2> XA4/CN0 0.06fF
C1884 XA3/XA4/MP2/a_216_n18# XA3/XA4/MP3/a_216_n18# 0.01fF
C1885 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128b<2>/XRES1A/B 0.03fF
C1886 XA5/DONE XA5/XA9/B 0.03fF
C1887 XA5/XA5/MN3/a_324_n18# XA5/CN0 0.01fF
C1888 XA6/XA1/XA1/MP3/G AVSS 0.13fF
C1889 XDAC1/XC1/XRES16/B SARP 21.64fF
C1890 XA3/XA3/MP2/a_216_n18# XA3/CN1 0.15fF
C1891 XA20/CNO XA2/XA1/XA1/MN2/S 0.03fF
C1892 XA3/XA8/MN0/a_324_n18# XA3/XA9/A 0.09fF
C1893 XA1/XA7/MP0/a_216_n18# AVDD 0.09fF
C1894 XA7/CN0 XA4/CN0 0.11fF
C1895 XB2/XA7/MN1/a_324_334# AVSS 0.08fF
C1896 XA7/XA1/XA5/MN2/S XA7/XA2/A 0.05fF
C1897 XA20/XA2/MP4/a_216_n18# XA20/XA9/Y 0.08fF
C1898 XA6/CP0 D<1> 0.01fF
C1899 D<2> XA5/CN0 0.06fF
C1900 XA20/XA3/N1 AVDD 1.01fF
C1901 XA8/ENO XA8/XA1/XA1/MP3/S 0.10fF
C1902 XA8/XA9/B XA8/XA9/MP1/a_216_n18# 0.07fF
C1903 XDAC2/XC64b<1>/XRES8/B XDAC2/XC0/XRES1A/B 0.03fF
C1904 XA8/XA1/XA4/MN2/S AVDD 0.02fF
C1905 XA4/XA1/XA2/Y XA20/CPO 0.22fF
C1906 XA1/XA12/MP0/a_216_n18# XA0/CEO 0.08fF
C1907 XB2/XA4/GNG XDAC2/XC1/XRES16/B 0.64fF
C1908 XA3/XA1/XA4/MN1/S XA3/EN 0.02fF
C1909 XDAC2/XC64b<1>/XRES1A/B XDAC2/XC64b<1>/XRES16/B 1.60fF
C1910 XA7/CN0 XA5/CN0 0.72fF
C1911 XA7/XA9/B XA8/XA9/B 0.07fF
C1912 D<3> XA4/CN0 0.12fF
C1913 XA7/XA9/MP1/a_216_n18# XA7/XA9/B 0.07fF
C1914 XA7/CEO VREF 0.04fF
C1915 XB2/XCAPB1/XCAPB3/m3_324_308# XB2/XA4/GNG 0.07fF
C1916 XDAC2/XC0/XRES2/B XDAC2/XC0/XRES8/B 1.58fF
C1917 XA0/XA1/XA5/MP1/S AVDD 0.13fF
C1918 XA6/CEO XA6/XA11/A 0.02fF
C1919 XA0/CP1 XDAC1/X16ab/XRES16/B 0.05fF
C1920 XB1/M4/G XA0/CEIN 0.26fF
C1921 XA2/XA2/MN2/a_324_n18# XA2/XA2/A 0.15fF
C1922 XDAC1/XC32a<0>/XRES4/B XDAC1/XC64a<0>/XRES4/B 0.10fF
C1923 XA5/XA2/MP2/a_216_n18# XA5/XA2/A 0.15fF
C1924 XA4/CN1 XA3/XA4/A 0.04fF
C1925 XA5/EN XA4/XA1/XA2/MN0/a_324_n18# 0.09fF
C1926 D<3> XA5/CN0 2.22fF
C1927 XA8/XA2/A XA8/XA4/A 0.14fF
C1928 XA8/CEO DONE 0.28fF
C1929 XA3/XA1/XA4/MP2/a_216_n18# XA3/XA1/XA4/MP1/a_216_n18# 0.01fF
C1930 XA5/CEO XA4/CEO 0.40fF
C1931 XA6/CN1 XA6/XA2/MN2/a_324_n18# 0.02fF
C1932 XA2/EN XA2/CN0 0.02fF
C1933 XA0/XA1/XA2/Y XA1/EN 0.10fF
C1934 XB2/XA3/B XB2/M4/G 0.06fF
C1935 XA2/CN0 XA2/XA6/MP2/a_216_n18# 0.08fF
C1936 XDAC1/XC64b<1>/XRES2/B SARP 3.05fF
C1937 XA5/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C1938 XA2/CN1 AVSS 2.46fF
C1939 XDAC1/XC1/XRES8/B XDAC1/XC64a<0>/XRES8/B 0.21fF
C1940 XA20/XA3a/A XA20/XA3a/MN0/a_324_n18# 0.08fF
C1941 XA7/XA9/Y AVDD 0.58fF
C1942 XA6/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C1943 CK_SAMPLE_BSSW XB1/XA3/MP0/a_216_n18# 0.08fF
C1944 XB2/M4/G AVSS 0.98fF
C1945 XA4/XA4/MP1/a_216_n18# XA4/XA4/MP0/a_216_n18# 0.01fF
C1946 VREF XA8/XA6/MP0/a_216_n18# 0.01fF
C1947 D<1> XA7/XA4/MP0/a_216_n18# 0.01fF
C1948 XB2/M4/G XB2/M5/a_324_n18# 0.07fF
C1949 XDAC2/XC1/XRES16/B XDAC2/XC64a<0>/XRES1A/B 0.04fF
C1950 XA20/XA3a/A XA20/XA3a/MN3/a_324_n18# 0.15fF
C1951 XA6/CN0 XA6/EN 0.03fF
C1952 XA20/XA11/MP0/a_216_n18# AVDD 0.09fF
C1953 XA3/XA5/MP1/a_216_n18# XA3/XA5/MP0/a_216_n18# 0.01fF
C1954 XA2/XA4/A XA2/XA3/MN3/a_324_n18# 0.01fF
C1955 AVDD XA20/XA9/MP0/a_216_n18# 0.17fF
C1956 XA20/XA1/MN1/a_324_n18# XA20/XA9/A 0.07fF
C1957 XA8/XA1/XA1/MP3/a_216_n18# XA20/CPO 0.08fF
C1958 XA20/XA1/MP0/S XA20/XA1/MN3/a_324_n18# 0.01fF
C1959 XA1/XA1/XA2/MN0/a_324_n18# XA1/XA1/XA1/MP3/G 0.06fF
C1960 XA0/CP0 XA0/CN0 4.08fF
C1961 XA2/XA2/A XA2/XA2/MN1/a_324_n18# 0.15fF
C1962 XA2/XA12/MP0/a_216_n18# XA2/XA11/MP1/a_216_n18# 0.01fF
C1963 AVDD XA0/CEIN 7.23fF
C1964 XA7/XA8/MP0/a_216_n18# AVDD 0.09fF
C1965 XA8/XA1/XA1/MN0/a_324_n18# AVSS 0.08fF
C1966 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MP3/S 0.04fF
C1967 XA0/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C1968 XA3/CP0 D<8> 0.03fF
C1969 XA8/XA5/MN0/a_324_n18# XA8/XA4/MN3/a_324_n18# 0.01fF
C1970 XA3/XA9/B XA3/XA6/MN1/S 0.05fF
C1971 XA4/XA11/A XA4/XA11/MN0/a_324_n18# 0.09fF
C1972 XA4/XA1/XA1/MN0/a_324_n18# XA4/XA1/XA1/MN1/a_324_n18# 0.01fF
C1973 XA20/XA13/MN1/a_324_334# AVSS 0.11fF
C1974 XA7/XA1/XA2/Y XA7/XA4/A 0.19fF
C1975 XA8/XA11/MP1/S AVDD 0.20fF
C1976 XA2/EN XA2/XA1/XA4/MN1/S 0.02fF
C1977 XA6/XA1/XA1/MP1/a_216_n18# XA6/XA1/XA1/MP3/G 0.01fF
C1978 XA6/XA1/XA2/Y XA6/EN 0.14fF
C1979 XA5/XA1/XA1/MP3/G AVSS 0.12fF
C1980 XA20/XA3a/A XA20/XA2/MP6/a_216_334# 0.01fF
C1981 XA5/XA1/XA4/MN2/S XA5/XA1/XA4/MP2/S 0.01fF
C1982 XA2/XA5/MN1/a_324_n18# XA2/XA5/MN0/a_324_n18# 0.01fF
C1983 XA4/XA1/XA1/MP1/a_216_n18# AVDD 0.08fF
C1984 XA5/CN0 XA5/XA5/MP3/a_216_n18# 0.02fF
C1985 D<3> XA5/XA6/MP3/a_216_n18# 0.15fF
C1986 D<2> XA6/CP0 0.23fF
C1987 XA2/XA4/MP0/a_216_n18# VREF 0.02fF
C1988 XA1/XA2/MP3/a_216_n18# XA1/CN1 0.02fF
C1989 XA3/XA2/MN2/a_324_n18# XA3/CN1 0.02fF
C1990 XA0/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C1991 XA7/XA9/B VREF 0.12fF
C1992 EN XA6/XA1/XA1/MP3/G 0.10fF
C1993 XA5/XA7/MP0/a_216_n18# D<3> 0.08fF
C1994 XA20/CPO XA6/XA1/XA1/MP3/a_216_n18# 0.08fF
C1995 XA7/XA11/A XA7/XA9/Y 0.14fF
C1996 XB2/XA3/MN0/a_324_n18# CK_SAMPLE_BSSW 0.07fF
C1997 XA4/XA4/MP0/a_216_n18# VREF 0.02fF
C1998 XA6/XA1/XA1/MP2/a_216_n18# XA6/XA1/XA1/MP3/a_216_n18# 0.01fF
C1999 XA20/XA1/MP2_DMY/a_216_n18# XA20/XA1/MP0/a_216_334# 0.01fF
C2000 XA7/XA3/MN2/a_324_n18# XA7/CN1 0.16fF
C2001 XDAC1/XC1/XRES1B/B XDAC1/XC1/XRES1A/B 0.01fF
C2002 XA0/XA9/MP1/a_216_334# AVDD 0.09fF
C2003 XA6/XA1/XA4/MP1/S XA7/EN 0.02fF
C2004 XA8/XA7/MP0/a_216_n18# AVDD 0.09fF
C2005 XA5/EN XA20/CPO 0.62fF
C2006 XA4/XA2/A XA4/XA2/MP0/a_216_n18# 0.08fF
C2007 XA3/EN XA2/XA1/XA2/Y 0.10fF
C2008 XDAC1/XC64b<1>/XRES16/B XDAC1/XC0/XRES16/B 0.41fF
C2009 XDAC2/XC128b<2>/XRES8/B AVSS 9.08fF
C2010 XA6/XA11/MN1/a_324_n18# AVSS 0.01fF
C2011 XA6/EN XA5/XA8/MN0/a_324_n18# 0.06fF
C2012 XA3/CN0 D<1> 0.04fF
C2013 XA20/XA3a/A XA20/XA3/MP0/a_216_n18# 0.09fF
C2014 XA1/XA11/MP1/a_216_n18# AVDD 0.08fF
C2015 XA5/XA4/A AVSS 1.11fF
C2016 XA6/XA2/A XA5/XA2/A 0.03fF
C2017 XDAC2/XC64b<1>/XRES1A/B SARN 1.50fF
C2018 XA0/XA1/XA5/MN1/S AVDD 0.02fF
C2019 D<7> XA1/XA6/MP3/S 0.02fF
C2020 D<7> AVSS 3.57fF
C2021 AVSS XA8/XA9/B 0.60fF
C2022 VREF XA2/XA11/A 0.02fF
C2023 XDAC2/XC128b<2>/XRES8/B XDAC2/XC128a<1>/XRES1B/B 0.02fF
C2024 XA0/CP0 XA0/XA5/MP3/a_216_n18# 0.15fF
C2025 AVDD XA2/XA1/XA1/MP3/S 0.14fF
C2026 XA1/CP0 AVDD 1.48fF
C2027 XA6/CN1 XA6/XA2/MP1/a_216_n18# 0.01fF
C2028 XA1/XA1/XA2/MP0/a_216_n18# XA1/XA1/XA4/MP0/a_216_n18# 0.01fF
C2029 XA2/CN1 EN 0.08fF
C2030 XA8/XA2/MP0/a_216_n18# EN 0.08fF
C2031 XA7/XA4/MN1/a_324_n18# XA7/CP0 0.03fF
C2032 XDAC1/XC128b<2>/XRES4/B XDAC1/XC128b<2>/XRES1A/B 0.29fF
C2033 XA4/XA1/XA5/MP2/a_216_n18# XA4/XA1/XA5/MP1/a_216_n18# 0.01fF
C2034 XDAC2/XC1/XRES8/B XDAC2/XC1/XRES2/B 1.58fF
C2035 XA4/XA1/XA5/MN2/S XA20/CNO 0.01fF
C2036 XA0/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C2037 XB1/XCAPB1/XCAPB4/m3_252_308# XB1/XA3/B 0.02fF
C2038 AVDD XA2/CEO 1.75fF
C2039 XA1/CP0 XDAC1/XC128b<2>/XRES16/B 0.01fF
C2040 XA8/XA11/MP0/a_216_n18# AVDD 0.09fF
C2041 XA8/XA3/MP3/a_216_n18# D<0> 0.02fF
C2042 XA7/XA1/XA1/MP2/S XA7/XA1/XA1/MP3/S 0.04fF
C2043 XA4/XA1/XA1/MN2/S AVSS 0.30fF
C2044 XA3/XA11/A XA3/XA11/MP1/a_216_n18# 0.08fF
C2045 XA3/XA2/MP0/a_216_n18# EN 0.08fF
C2046 XA0/XA2/MN3/a_324_n18# D<8> 0.03fF
C2047 XA1/XA4/A XA0/XA4/A 0.03fF
C2048 XA1/EN XA0/XA1/XA1/MN2/S 0.06fF
C2049 CK_SAMPLE XA8/XA6/MN3/a_324_n18# 0.15fF
C2050 XDAC1/XC128b<2>/XRES8/B XDAC1/X16ab/XRES1A/B 0.03fF
C2051 XA7/XA4/MP1/a_216_n18# XA7/CP0 0.02fF
C2052 XA3/XA9/Y XA2/CEO 0.03fF
C2053 XA7/XA6/MN2/a_324_n18# AVSS 0.01fF
C2054 XA7/XA1/XA1/MN0/a_324_n18# XA7/EN 0.09fF
C2055 XA6/XA1/XA4/MN1/a_324_n18# XA6/XA1/XA4/MN2/a_324_n18# 0.01fF
C2056 XA3/XA11/MP1/S XA3/XA12/A 0.06fF
C2057 XA7/CN1 XA7/EN 0.04fF
C2058 AVDD XA20/XA3a/MP0/a_216_n18# 0.09fF
C2059 XA2/XA3/MN1/a_324_n18# D<6> 0.02fF
C2060 XB2/XA4/GNG XB2/XA5/MP1/a_216_334# 0.01fF
C2061 XA5/XA1/XA1/MP3/G EN 0.10fF
C2062 XA0/XA1/XA5/MP2/S XA0/XA1/XA5/MN2/S 0.01fF
C2063 XA3/CN0 XA3/CN1 2.64fF
C2064 XA0/CP0 D<6> 0.22fF
C2065 XA7/XA9/MN1/a_324_334# XA7/XA9/MN1/a_324_n18# 0.01fF
C2066 D<7> XA1/XA3/MN1/a_324_n18# 0.02fF
C2067 XDAC1/XC0/XRES8/B XDAC1/XC0/XRES16/B 1.42fF
C2068 XA6/XA1/XA5/MP2/S AVDD 0.08fF
C2069 XA0/CP0 XA0/XA4/A 0.57fF
C2070 XB2/XA5b/MN1/a_324_n18# AVSS 0.12fF
C2071 XA2/CN1 XA2/XA2/MP1/a_216_n18# 0.02fF
C2072 XA7/XA1/XA5/MN1/a_324_n18# XA7/XA1/XA5/MN0/a_324_n18# 0.01fF
C2073 XA7/XA9/A XA7/XA9/MN0/a_324_n18# 0.15fF
C2074 XA6/CP0 XA8/EN 0.03fF
C2075 XA2/XA6/MN0/a_324_n18# XA2/XA5/MN3/a_324_n18# 0.01fF
C2076 XA3/XA1/XA1/MN3/a_324_n18# XA3/XA1/XA2/MN0/a_324_n18# 0.01fF
C2077 XA1/XA6/MP3/S VREF 0.02fF
C2078 XA20/XA12/Y VREF 0.03fF
C2079 VREF AVSS 8.49fF
C2080 XB2/XA1/MP0/G AVSS 0.21fF
C2081 XA5/XA1/XA2/MP0/a_216_n18# XA5/XA1/XA4/MP0/a_216_n18# 0.01fF
C2082 XA20/CNO XA2/XA1/XA1/MP2/a_216_n18# 0.08fF
C2083 D<7> CK_SAMPLE 0.10fF
C2084 CK_SAMPLE XA8/XA9/B 0.12fF
C2085 XA2/XA11/MP0/a_216_n18# XA2/XA9/MP1/a_216_334# 0.01fF
C2086 XB2/M4/G XB2/XA4/MN1/a_324_n18# 0.01fF
C2087 XA8/XA6/MP0/a_216_n18# XA8/CP0 0.08fF
C2088 XDAC1/XC64b<1>/XRES1A/B XDAC1/X16ab/XRES8/B 0.03fF
C2089 D<2> XA3/CN0 0.06fF
C2090 XA7/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C2091 XB1/XA3/MP0/S XB1/XA3/B 0.11fF
C2092 XDAC1/XC32a<0>/XRES8/B XDAC1/XC128a<1>/XRES16/B 0.03fF
C2093 XA2/XA11/MN0/a_324_n18# XA2/XA11/MN1/a_324_n18# 0.01fF
C2094 XA0/CEIN XB1/M6/a_324_n18# 0.15fF
C2095 XA5/XA1/XA1/MP3/G XA5/XA1/XA2/MN0/a_324_n18# 0.06fF
C2096 D<0> DONE 0.01fF
C2097 XA6/XA9/B XA6/XA12/A 0.01fF
C2098 XDAC1/X16ab/XRES4/B SARP 6.32fF
C2099 XDAC2/X16ab/XRES1B/B XDAC2/X16ab/XRES8/B 0.12fF
C2100 XA4/XA1/XA1/MP3/S XA4/XA1/XA1/MP2/S 0.04fF
C2101 XA7/XA5/MP2/a_216_n18# XA7/CP0 0.15fF
C2102 XA20/XA2/MP3/a_216_n18# XA20/XA2/MP2/a_216_n18# 0.01fF
C2103 XA4/XA1/XA1/MP1/a_216_n18# XA5/EN 0.01fF
C2104 XA5/XA6/MP2/a_216_n18# AVDD 0.09fF
C2105 XA3/CN0 XA7/CN0 0.09fF
C2106 XA1/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C2107 XA5/XA4/A EN 0.09fF
C2108 XDAC1/XC1/XRES1A/B SARP 1.51fF
C2109 XA3/XA1/XA1/MP1/a_216_n18# XA3/XA1/XA1/MP3/G 0.01fF
C2110 XDAC2/XC128a<1>/XRES1A/B SARN 1.50fF
C2111 XA4/XA1/XA4/MP1/S AVDD 0.14fF
C2112 CK_SAMPLE XA8/XA6/MP3/S 0.01fF
C2113 D<7> EN 0.05fF
C2114 XA20/XA2/MN0/a_324_n18# XA20/XA1/MN6/a_324_n18# 0.01fF
C2115 XA5/XA9/B VREF 0.12fF
C2116 XA7/XA3/MP2/a_216_n18# XA7/XA3/MP3/a_216_n18# 0.01fF
C2117 XA7/XA3/MP1/a_216_n18# XA7/CN1 0.15fF
C2118 XB1/XA1/MP0/G XB1/XA4/GNG 0.06fF
C2119 XA2/XA9/B VREF 0.12fF
C2120 XA3/XA1/XA1/MP3/G XA3/XA1/XA2/MN0/a_324_n18# 0.06fF
C2121 XA3/CN0 D<3> 0.11fF
C2122 XA0/XA1/XA4/MP2/S AVDD 0.11fF
C2123 XA1/XA1/XA2/Y XA1/EN 0.14fF
C2124 XA20/XA2/N2 XA20/CNO 0.04fF
C2125 XA5/XA6/MP0/a_216_n18# XA5/CN0 0.08fF
C2126 XA0/CP0 SARP 0.80fF
C2127 XA1/XA11/MN0/a_324_n18# XA1/XA9/MN1/a_324_334# 0.01fF
C2128 XA3/XA11/MP0/a_216_n18# XA3/XA11/A 0.07fF
C2129 XA0/CP1 XA3/CP0 0.06fF
C2130 XA4/EN XA2/XA1/XA1/MP3/G 0.01fF
C2131 XA8/CEO XA20/XA13/MP1/a_216_n18# 0.08fF
C2132 D<5> XA3/XA9/A 0.01fF
C2133 XA6/XA9/Y VREF 0.03fF
C2134 XA4/XA1/XA2/Y XA4/XA1/XA4/MP1/S 0.01fF
C2135 XA2/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C2136 XA7/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C2137 XA0/XA1/XA4/MP0/a_216_n18# XA0/XA1/XA2/MP0/a_216_n18# 0.01fF
C2138 XA20/XA13/MP1/a_216_334# AVSS 0.02fF
C2139 XB2/XA4/GNG XB2/XCAPB1/XCAPB2/m3_252_308# 0.13fF
C2140 XA8/XA9/A XA8/XA9/MP1/a_216_n18# 0.08fF
C2141 XA8/XA6/MN3/S XA8/XA9/B 0.09fF
C2142 XA8/XA1/XA2/Y AVSS 0.32fF
C2143 XA2/XA6/MP3/a_216_n18# XA2/XA6/MP2/a_216_n18# 0.01fF
C2144 XA2/XA9/MN1/a_324_n18# XA2/XA9/MN1/a_324_334# 0.01fF
C2145 XA5/CP0 XA5/XA5/MN3/a_324_n18# 0.15fF
C2146 XA0/CP0 XA0/XA5/MN0/a_324_n18# 0.09fF
C2147 XA1/XA4/A XA1/XA4/MP0/a_216_n18# 0.07fF
C2148 XA4/XA5/MN0/a_324_n18# XA4/XA4/MN3/a_324_n18# 0.01fF
C2149 XA7/XA9/B XA8/XA9/A 0.02fF
C2150 XDAC2/XC128b<2>/XRES16/B XDAC2/X16ab/XRES1A/B 0.04fF
C2151 XA5/XA1/XA1/MP2/S XA6/EN 0.14fF
C2152 XA20/CNO XA20/XA3a/A 0.24fF
C2153 XA20/XA13/MN1/a_324_n18# XA20/XA12/MN0/a_324_n18# 0.01fF
C2154 XA2/CN0 XA2/XA1/XA1/MP3/G 0.02fF
C2155 XA1/XA3/MP2/a_216_n18# XA1/CN1 0.15fF
C2156 XA7/XA6/MP1/a_216_n18# AVDD 0.08fF
C2157 VREF CK_SAMPLE 1.85fF
C2158 XDAC2/XC0/XRES16/B XDAC2/XC0/XRES4/B 0.25fF
C2159 AVDD XA2/XA1/XA0/MP1/a_216_n18# 0.15fF
C2160 XA6/XA6/MP1/a_216_n18# XA6/CN0 0.15fF
C2161 XDAC2/XC64a<0>/XRES16/B XDAC2/XC64a<0>/XRES2/B 1.61fF
C2162 XA0/XA1/XA4/MN2/S XA0/XA1/XA2/Y 0.05fF
C2163 XA1/XA11/MP0/a_216_n18# AVDD 0.09fF
C2164 XA7/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C2165 XA0/XA1/XA1/MP3/G XA1/EN 0.27fF
C2166 D<1> XA20/CNO 0.06fF
C2167 AVDD XA2/XA1/XA5/MP1/S 0.13fF
C2168 XA5/XA9/MN0/a_324_n18# XA5/XA9/A 0.15fF
C2169 XA7/XA2/MP3/a_216_n18# VREF 0.03fF
C2170 XA6/XA7/MN0/a_324_n18# XA6/XA8/MN0/a_324_n18# 0.01fF
C2171 XB2/XA5b/MN1/a_324_n18# XB2/XA0/MN0/a_324_n18# 0.01fF
C2172 XA3/XA2/MN2/a_324_n18# XA3/XA2/MN1/a_324_n18# 0.01fF
C2173 XB1/XA4/MN1/a_324_n18# XB1/XA1/Y 0.08fF
C2174 AVDD XA8/XA9/Y 0.59fF
C2175 XDAC1/XC0/XRES1B/B SARP 1.84fF
C2176 XA20/XA2/MP4/a_216_n18# AVDD 0.09fF
C2177 XA1/XA9/B XA1/XA6/MN1/S 0.05fF
C2178 XA8/XA5/MP2/a_216_n18# XA8/XA5/MP3/a_216_n18# 0.01fF
C2179 EN VREF 1.75fF
C2180 XA6/EN XA5/XA1/XA1/MP3/a_216_n18# 0.01fF
C2181 XA5/XA7/MN0/a_324_n18# XA5/XA8/MN0/a_324_n18# 0.01fF
C2182 XA20/XA4/MP2_DMY/a_216_n18# XA20/XA4/MP0/a_216_334# 0.01fF
C2183 XB1/CKN XB1/XA4/MN1/a_324_n18# 0.07fF
C2184 XA7/XA9/A AVDD 0.62fF
C2185 XA20/XA4/MP0/S AVSS 0.45fF
C2186 EN XA0/XA1/XA5/MN0/a_324_n18# 0.07fF
C2187 XA0/XA2/MN2/a_324_n18# XA0/XA2/MN1/a_324_n18# 0.01fF
C2188 XA5/CP0 D<3> 0.23fF
C2189 D<3> XA5/XA6/MP1/a_216_n18# 0.01fF
C2190 XA20/XA10/MN1/S XA20/XA9/A 0.13fF
C2191 AVDD XA0/XA6/MN1/S 0.01fF
C2192 XA1/EN D<8> 0.12fF
C2193 XA8/EN XA7/XA1/XA5/MP1/S 0.02fF
C2194 XA4/EN XA3/XA4/A 0.12fF
C2195 XA6/XA1/XA4/MN2/a_324_n18# XA6/EN 0.08fF
C2196 XA2/XA4/A XA2/XA1/XA5/MP2/S 0.02fF
C2197 XDAC1/XC32a<0>/XRES4/B XDAC1/XC128a<1>/XRES1A/B 0.01fF
C2198 XA5/XA3/MN2/a_324_n18# XA5/CN1 0.16fF
C2199 XDAC1/XC128b<2>/XRES1A/B AVSS 2.95fF
C2200 XA1/XA3/MP1/a_216_n18# XA1/CN1 0.15fF
C2201 D<0> XA8/XA6/MN1/S 0.01fF
C2202 XA3/XA6/MP3/a_216_n18# XA3/XA7/MP0/a_216_n18# 0.01fF
C2203 XA3/XA9/B XA3/XA9/MN1/a_324_n18# 0.09fF
C2204 VREF XA2/XA12/A 0.03fF
C2205 XA3/XA5/MP1/a_216_n18# AVDD 0.07fF
C2206 XA20/XA9/Y XA20/XA2/MP2/a_216_n18# 0.08fF
C2207 XA7/CEO XA8/XA11/MN1/a_324_n18# 0.08fF
C2208 XA20/XA3/N2 AVSS 0.23fF
C2209 XDAC2/XC1/XRES2/B XDAC2/XC64a<0>/XRES16/B 0.01fF
C2210 XA7/XA9/MN1/a_324_334# XA7/XA9/Y 0.09fF
C2211 XA2/XA8/MP0/a_216_n18# AVDD 0.09fF
C2212 XA7/CN0 XA7/XA5/MN3/a_324_n18# 0.01fF
C2213 XA3/XA1/XA1/MP3/a_216_n18# XA3/XA1/XA1/MP3/G 0.07fF
C2214 XA4/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C2215 XA2/XA9/A XA3/EN 0.09fF
C2216 XA3/XA2/A AVSS 0.24fF
C2217 XA8/XA9/B XA8/XA9/MN1/S 0.02fF
C2218 XDAC1/XC128a<1>/XRES1A/B XDAC1/XC128a<1>/XRES4/B 0.29fF
C2219 XDAC1/XC128a<1>/XRES2/B XDAC1/XC128a<1>/XRES1B/B 0.23fF
C2220 XDAC1/XC1/XRES8/B XDAC1/XC1/XRES4/B 2.60fF
C2221 XA1/XA6/MN3/a_324_n18# XA1/XA7/MN0/a_324_n18# 0.01fF
C2222 VREF XA2/XA2/MP1/a_216_n18# 0.02fF
C2223 XA5/XA9/A XA5/XA8/MP0/a_216_n18# 0.07fF
C2224 XA8/XA1/XA1/MP1/a_216_n18# XA8/XA1/XA1/MP2/a_216_n18# 0.01fF
C2225 XA3/XA6/MN1/S AVSS 0.15fF
C2226 XA7/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C2227 XA4/XA2/MP1/a_216_n18# AVDD 0.08fF
C2228 XA7/XA11/MN1/a_324_n18# XA6/CEO 0.08fF
C2229 XA8/ENO DONE 0.06fF
C2230 XB1/XCAPB1/XCAPB1/m3_9828_132# XB1/XA4/GNG 0.04fF
C2231 AVSS XA8/CP0 0.92fF
C2232 XA5/EN XA4/XA1/XA4/MP1/S 0.02fF
C2233 XA3/XA2/A XA3/XA2/MN3/a_324_n18# 0.15fF
C2234 XA20/CNO XA3/CN1 0.23fF
C2235 XA6/CN0 XA2/CN0 0.05fF
C2236 XB2/XA3/MP0/S CK_SAMPLE_BSSW 0.01fF
C2237 XA1/XA1/XA4/MN2/S XA20/CNO 0.01fF
C2238 XA7/XA11/A XA7/XA9/A 0.01fF
C2239 XA7/XA2/MP1/a_216_n18# XA7/XA2/MP0/a_216_n18# 0.01fF
C2240 XA6/XA8/MP0/a_216_n18# XA7/EN 0.08fF
C2241 XDAC2/XC1/XRES4/B XDAC2/XC1/XRES16/B 0.25fF
C2242 XA7/XA1/XA1/MP3/G AVDD 0.62fF
C2243 XA8/XA1/XA2/Y EN 0.06fF
C2244 XA3/XA1/XA1/MP2/S AVDD 0.09fF
C2245 XA5/CP0 XA5/XA5/MP3/a_216_n18# 0.15fF
C2246 XDAC2/XC32a<0>/XRES4/B AVSS 5.78fF
C2247 SARP CK_SAMPLE_BSSW 0.01fF
C2248 XA8/EN XA7/XA7/MN0/a_324_n18# 0.08fF
C2249 XA4/XA9/A VREF 0.04fF
C2250 XA2/XA3/MN0/a_324_n18# XA2/XA2/A 0.07fF
C2251 XA7/XA1/XA2/Y XA7/EN 0.14fF
C2252 XDAC1/XC0/XRES8/B XA1/CN1 0.02fF
C2253 XA8/CN1 VREF 0.70fF
C2254 XDAC2/XC128a<1>/XRES8/B XDAC2/XC32a<0>/XRES8/B 0.21fF
C2255 XA20/CPO XA1/CN1 0.19fF
C2256 XA6/CN1 XA6/XA3/MN1/a_324_n18# 0.16fF
C2257 XB2/M6/a_324_n18# SARP 0.01fF
C2258 AVDD XA2/XA13/MP1/a_216_334# 0.17fF
C2259 D<2> XA20/CNO 0.06fF
C2260 XDAC2/XC64a<0>/XRES8/B AVSS 9.11fF
C2261 XA8/XA9/A AVSS 0.31fF
C2262 XA8/XA2/MP2/a_216_n18# AVDD 0.07fF
C2263 XA7/XA2/MP1/a_216_n18# XA7/CN1 0.01fF
C2264 XA6/XA6/MN3/S AVDD 0.01fF
C2265 AVDD XA2/XA1/XA5/MN1/S 0.02fF
C2266 XA7/XA5/MN0/a_324_n18# XA7/XA4/A 0.07fF
C2267 XA4/XA2/MN3/a_324_n18# XA4/XA3/MN0/a_324_n18# 0.01fF
C2268 CK_SAMPLE XA20/XA4/MP0/S 0.06fF
C2269 XA1/CP0 XA1/XA2/A 0.04fF
C2270 XB1/M2/a_324_n18# XB1/M3/a_324_n18# 0.01fF
C2271 XA7/CN0 XA20/CNO 0.06fF
C2272 XA1/XA4/A XA1/XA4/MN1/a_324_n18# 0.15fF
C2273 XA6/CN0 SARN 0.07fF
C2274 XA4/XA11/MP1/a_216_n18# AVDD 0.08fF
C2275 XA3/XA3/MN0/a_324_n18# XA3/XA2/MN3/a_324_n18# 0.01fF
C2276 XA1/CEO XA1/XA11/MP1/S 0.02fF
C2277 XA6/XA2/A XA7/EN 0.10fF
C2278 XA8/XA1/XA4/MP1/a_216_n18# XA8/XA1/XA4/MP2/a_216_n18# 0.01fF
C2279 XA0/XA3/MP1/a_216_n18# XA0/XA3/MP2/a_216_n18# 0.01fF
C2280 XA5/XA12/A XA5/XA12/MP0/a_216_n18# 0.07fF
C2281 XA0/XA12/A AVDD 0.44fF
C2282 XA0/XA1/XA2/Y XA0/CN0 0.02fF
C2283 XDAC2/XC0/XRES1B/B XDAC2/XC0/XRES4/B 1.64fF
C2284 D<1> XA7/XA3/MP2/a_216_n18# 0.01fF
C2285 D<3> XA20/CNO 0.06fF
C2286 XA3/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C2287 XA4/XA1/XA1/MP3/a_216_n18# XA20/CPO 0.08fF
C2288 XA7/XA9/B XA7/XA9/MN1/a_324_n18# 0.09fF
C2289 XA4/XA2/A AVSS 0.26fF
C2290 XA0/XA4/A XA0/XA5/MP0/a_216_n18# 0.08fF
C2291 XB2/XA1/Y AVDD 0.45fF
C2292 XA4/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C2293 XA20/XA4/MP5_DMY/a_216_n18# XA20/XA4/MP4_DMY/a_216_n18# 0.01fF
C2294 XA7/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C2295 XA0/XA6/MP3/S XA0/XA9/B 0.07fF
C2296 XA6/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C2297 XA5/XA1/XA1/MP0/a_216_n18# AVDD 0.14fF
C2298 XA20/XA9/A XA20/XA4/MP0/a_216_n18# 0.06fF
C2299 XA3/CP0 XA4/EN 0.14fF
C2300 XA2/XA4/A XA2/XA2/A 0.14fF
C2301 XA8/XA11/MN1/a_324_n18# XA8/XA11/MN0/a_324_n18# 0.01fF
C2302 XA1/XA1/XA4/MN1/a_324_n18# XA1/XA1/XA4/MN0/a_324_n18# 0.01fF
C2303 XDAC1/XC1/XRES16/B XB1/XA4/GNG 0.65fF
C2304 XA7/XA1/XA5/MN2/S AVSS 0.09fF
C2305 XA3/XA6/MN1/S CK_SAMPLE 0.05fF
C2306 XA6/XA9/B XA6/XA9/MP1/a_216_334# 0.08fF
C2307 XA7/XA1/XA1/MN2/S XA20/CNO 0.03fF
C2308 CK_SAMPLE XA8/CP0 0.08fF
C2309 XB2/XA7/MN1/a_324_n18# AVSS 0.09fF
C2310 XB2/XA4/GNG XB2/XA3/MP0/S 0.02fF
C2311 XA8/EN XA7/XA1/XA4/MP2/S 0.02fF
C2312 XA6/XA9/MN1/S AVDD 0.01fF
C2313 XA5/CN0 XA5/XA6/MP1/S 0.02fF
C2314 XA3/XA3/MP0/a_216_n18# XA3/CN1 0.07fF
C2315 XA1/XA8/MP0/a_216_n18# XA1/XA7/MP0/a_216_n18# 0.01fF
C2316 XA4/XA13/MN1/a_324_n18# AVSS 0.09fF
C2317 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128a<1>/XRES8/B 0.03fF
C2318 XA3/XA2/A EN 0.11fF
C2319 XA4/XA9/B XA4/XA12/A 0.01fF
C2320 XA5/XA5/MP0/a_216_n18# XA5/XA4/A 0.08fF
C2321 VREF XA2/XA4/MP3/a_216_n18# 0.03fF
C2322 XA8/XA3/MP2/a_216_n18# XA8/XA3/MP1/a_216_n18# 0.01fF
C2323 XA8/EN XA7/XA1/XA4/MN0/a_324_n18# 0.07fF
C2324 XA0/CEIN XB1/XA1/Y 0.07fF
C2325 XA4/XA2/MN3/a_324_n18# XA4/XA2/MN2/a_324_n18# 0.01fF
C2326 XA7/XA1/XA4/MN1/S AVSS 0.10fF
C2327 XA6/XA9/MP1/a_216_n18# XA6/XA9/MP1/a_216_334# 0.01fF
C2328 XA20/CPO XA3/XA1/XA1/MP3/G 0.15fF
C2329 XA7/XA4/MP0/a_216_n18# XA7/CN1 0.08fF
C2330 XA7/XA1/XA4/MN2/S XA7/XA4/A 0.06fF
C2331 XA2/CN0 XA3/CP0 0.04fF
C2332 XA5/XA3/MP0/a_216_n18# VREF 0.02fF
C2333 XA5/XA1/XA1/MN1/a_324_n18# XA5/EN 0.07fF
C2334 XA2/XA9/Y XA2/XA9/A 0.04fF
C2335 XA0/CEIN XB1/CKN 0.08fF
C2336 XA1/XA1/XA1/MP3/S AVSS 0.02fF
C2337 XA6/XA9/B AVDD 0.79fF
C2338 XA6/XA1/XA4/MN2/S AVSS 0.06fF
C2339 XA5/XA9/Y XA5/XA9/MP1/a_216_334# 0.07fF
C2340 CK_SAMPLE XA8/XA9/A 0.05fF
C2341 XB1/XA3/MP0/S XB1/XA3/MN1/a_324_n18# 0.01fF
C2342 XA4/XA2/MP2/a_216_n18# VREF 0.03fF
C2343 SAR_IN XB2/XA3/MP0/S 0.06fF
C2344 XA0/XA1/XA1/MP3/S AVSS 0.02fF
C2345 XA6/EN XA5/XA1/XA2/Y 0.14fF
C2346 XA6/XA1/XA4/MN1/S XA6/EN 0.02fF
C2347 D<5> XDAC1/X16ab/XRES16/B 0.07fF
C2348 XA6/CN0 XA6/XA4/A 0.12fF
C2349 XB2/XA2/MP0/G AVSS 0.09fF
C2350 XA8/EN XA8/XA1/XA5/MN0/a_324_n18# 0.07fF
C2351 SAR_IN SARP 0.59fF
C2352 XA6/XA2/MP1/a_216_n18# XA6/XA2/MP0/a_216_n18# 0.01fF
C2353 D<7> XA2/CN1 0.09fF
C2354 XA6/XA9/MP1/a_216_n18# AVDD 0.09fF
C2355 XDAC1/XC128a<1>/XRES2/B XDAC1/XC128b<2>/XRES16/B 0.01fF
C2356 XA3/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C2357 XA3/XA9/A AVDD 0.62fF
C2358 XA4/XA3/MN1/a_324_n18# XA4/CN1 0.16fF
C2359 XA4/XA11/MP1/a_216_n18# XA4/XA12/MP0/a_216_n18# 0.01fF
C2360 XB1/XA4/GNG XB1/XA7/MP1/a_216_n18# 0.02fF
C2361 XA3/CP0 SARN 0.03fF
C2362 XA8/EN XA20/CNO 0.99fF
C2363 XA5/XA1/XA1/MP0/a_216_n18# XA5/XA1/XA0/MP1/a_216_n18# 0.01fF
C2364 XA0/XA2/A AVDD 1.07fF
C2365 XA3/XA5/MP3/a_216_n18# XA3/XA6/MP0/a_216_n18# 0.01fF
C2366 XA0/CP1 XA1/EN 0.42fF
C2367 XA2/CP0 D<4> 0.26fF
C2368 XA6/XA1/XA2/Y XA6/XA4/A 0.19fF
C2369 XA1/XA1/XA1/MP2/a_216_n18# XA20/CNO 0.08fF
C2370 XA4/CN0 XA4/XA4/A 0.12fF
C2371 XA3/XA9/Y XA3/XA9/A 0.04fF
C2372 XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MP1/a_216_n18# 0.01fF
C2373 XA0/XA1/XA2/Y XA0/XA1/XA4/MP1/S 0.01fF
C2374 XA7/CEO XA7/XA9/Y 0.04fF
C2375 XB1/XCAPB1/XCAPB1/m3_324_308# XB1/XA4/GNG 0.07fF
C2376 XA0/XA2/A XA0/XA2/MP1/a_216_n18# 0.15fF
C2377 XA2/EN AVDD 4.10fF
C2378 XA4/XA9/B XA4/XA11/A 0.03fF
C2379 XA2/XA6/MP2/a_216_n18# AVDD 0.09fF
C2380 XA3/XA9/B XA2/CEO 0.02fF
C2381 XA7/XA1/XA4/MP1/S AVDD 0.14fF
C2382 XA6/XA4/MN2/a_324_n18# AVSS 0.01fF
C2383 XA1/XA6/MP3/a_216_n18# AVDD 0.08fF
C2384 XA5/XA1/XA1/MN1/a_324_n18# XA5/XA1/XA1/MN0/a_324_n18# 0.01fF
C2385 XDAC2/XC128b<2>/XRES16/B D<8> 0.05fF
C2386 XA8/XA11/MN1/a_324_n18# AVSS 0.01fF
C2387 XA4/XA2/A EN 0.14fF
C2388 XA1/XA1/XA2/Y XA1/XA1/XA4/MN0/a_324_n18# 0.02fF
C2389 XA1/CEO XA0/CEO 0.41fF
C2390 XA8/XA4/MN0/a_324_n18# XA8/XA3/MN3/a_324_n18# 0.01fF
C2391 XA6/XA9/A D<2> 0.01fF
C2392 XA5/CP0 XA5/XA6/MP0/a_216_n18# 0.08fF
C2393 XA5/XA6/MP0/a_216_n18# XA5/XA6/MP1/a_216_n18# 0.01fF
C2394 XA8/CN1 XA8/CP0 0.03fF
C2395 XA4/XA4/A XA4/XA4/MN0/a_324_n18# 0.09fF
C2396 XA5/XA5/MP0/a_216_n18# VREF 0.02fF
C2397 XA7/XA1/XA5/MN2/S EN 0.02fF
C2398 XA0/XA1/XA4/MN1/a_324_n18# XA0/XA1/XA4/MN0/a_324_n18# 0.01fF
C2399 XDAC2/XC128a<1>/XRES16/B D<8> 0.22fF
C2400 D<3> XA5/XA9/A 0.01fF
C2401 XA0/XA4/A XA0/XA1/XA2/Y 0.19fF
C2402 XA0/XA9/MP1/a_216_n18# XA0/XA9/B 0.07fF
C2403 XA0/XA6/MP3/a_216_n18# XA0/XA6/MP2/a_216_n18# 0.01fF
C2404 XDAC1/XC64b<1>/XRES16/B AVSS 16.03fF
C2405 XB2/M2/a_324_n18# XB2/M4/G 0.15fF
C2406 XA1/XA1/XA4/MN1/S AVSS 0.10fF
C2407 XDAC2/X16ab/XRES1A/B XDAC2/X16ab/XRES2/B 0.25fF
C2408 XA3/XA1/XA5/MP1/a_216_n18# XA3/XA1/XA5/MP0/a_216_n18# 0.01fF
C2409 XA1/CP0 XA1/CN1 0.20fF
C2410 XA7/XA1/XA5/MN2/a_324_n18# XA7/EN 0.08fF
C2411 XDAC2/XC128a<1>/XRES4/B XDAC2/XC128a<1>/XRES8/B 2.60fF
C2412 XDAC2/XC64b<1>/XRES1A/B XDAC2/XC64b<1>/XRES2/B 0.25fF
C2413 XA7/XA1/XA1/MP3/S XA20/CPO 0.01fF
C2414 XA7/XA1/XA4/MP0/a_216_n18# XA7/XA1/XA2/MP0/a_216_n18# 0.01fF
C2415 XA3/XA13/MN1/a_324_n18# XA3/XA13/MN1/a_324_334# 0.01fF
C2416 EN XA0/XA1/XA4/MP0/a_216_n18# 0.07fF
C2417 XA3/XA5/MP0/a_216_n18# XA3/XA4/A 0.08fF
C2418 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC64a<0>/XRES1B/B 0.03fF
C2419 XDAC1/X16ab/XRES4/B XDAC1/X16ab/XRES8/B 2.60fF
C2420 XA8/XA1/XA4/MP1/a_216_n18# XA8/XA1/XA4/MP0/a_216_n18# 0.01fF
C2421 XA20/XA4/MN5/a_324_n18# XA20/XA4/MP0/S 0.01fF
C2422 XA0/XA12/MP0/a_216_n18# XA0/CEIN 0.08fF
C2423 XA7/XA1/XA1/MP3/G XA7/XA1/XA2/MP0/a_216_n18# 0.08fF
C2424 XDAC1/XC32a<0>/XRES16/B AVSS 17.65fF
C2425 XB1/XA3/MP0/S XB1/XA4/MN0/a_324_n18# 0.07fF
C2426 XDAC1/XC64b<1>/XRES16/B XDAC1/X16ab/XRES1B/B 0.05fF
C2427 XA0/XA5/MN1/a_324_n18# XA0/CN0 0.02fF
C2428 XB2/XA4/MN1/a_324_334# AVSS 0.01fF
C2429 XA1/XA1/XA2/MP0/a_216_n18# XA1/XA1/XA1/MP3/G 0.08fF
C2430 XA2/XA9/MN1/a_324_n18# XA2/XA9/B 0.09fF
C2431 XA0/XA11/MN1/a_324_n18# AVSS 0.01fF
C2432 XA0/CP0 XA0/XA4/MP3/a_216_n18# 0.02fF
C2433 XDAC1/XC128b<2>/XRES1A/B XDAC1/X16ab/XRES1A/B 0.03fF
C2434 XA1/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C2435 D<0> XA20/CNO 0.01fF
C2436 XA2/CN1 VREF 0.77fF
C2437 XA5/XA1/XA1/MP0/a_216_n18# XA5/EN 0.01fF
C2438 AVDD XA8/XA5/MP2/a_216_n18# 0.07fF
C2439 XA2/XA1/XA5/MN2/S XA2/XA1/XA5/MP2/S 0.01fF
C2440 XA4/XA5/MP0/a_216_n18# VREF 0.02fF
C2441 XA4/XA3/MN2/a_324_n18# XA4/XA4/A 0.01fF
C2442 XA6/XA1/XA2/MP0/a_216_n18# XA7/EN 0.08fF
C2443 XA4/XA2/MN2/a_324_n18# XA4/XA2/MN1/a_324_n18# 0.01fF
C2444 XB2/M4/G XB2/XA1/MP0/G 0.04fF
C2445 XA5/XA4/MN0/a_324_n18# XA5/XA3/MN3/a_324_n18# 0.01fF
C2446 XA1/XA1/XA1/MN1/a_324_n18# XA1/EN 0.07fF
C2447 XA0/XA9/Y AVSS 0.21fF
C2448 XA20/XA1/MN5/a_324_n18# XA20/XA1/MP0/S 0.01fF
C2449 XA20/XA9/MP0/a_216_334# XA20/XA9/MP0/a_216_n18# 0.01fF
C2450 XA4/XA5/MN1/a_324_n18# XA4/CN0 0.02fF
C2451 XA7/XA9/B XA7/XA9/Y 0.15fF
C2452 XB1/XA0/MP0/a_216_n18# XB1/XA3/B 0.01fF
C2453 XA4/XA6/MP0/a_216_n18# XA4/CP0 0.08fF
C2454 XB2/CKN XB2/XA3/B 0.29fF
C2455 XA3/XA3/MN2/a_324_n18# XA3/XA3/MN1/a_324_n18# 0.01fF
C2456 XB2/XA4/GNG XB2/XCAPB1/XCAPB4/m3_9756_132# 0.02fF
C2457 XA4/XA6/MP1/S AVDD 0.12fF
C2458 XA20/XA10/MN1/S AVDD 0.01fF
C2459 XA0/XA4/MP2/a_216_n18# AVDD 0.07fF
C2460 XA1/XA9/B XA1/CN0 0.07fF
C2461 XA20/XA2/MN4/a_324_n18# XA20/XA2/MN3/a_324_n18# 0.01fF
C2462 XA8/XA6/MP3/S XA8/XA9/B 0.07fF
C2463 XA1/XA1/XA1/MN2/S AVDD 0.05fF
C2464 XDAC1/XC128b<2>/XRES8/B XDAC1/XC128b<2>/XRES1A/B 0.12fF
C2465 D<5> XA3/XA4/A 0.26fF
C2466 XA20/XA2/MP6/a_216_n18# AVDD 0.09fF
C2467 XB2/CKN AVSS 0.71fF
C2468 XA20/CPO XA0/XA1/XA4/MN0/a_324_n18# 0.09fF
C2469 XA1/XA6/MP2/a_216_n18# XA1/CN0 0.08fF
C2470 XA6/XA9/Y XA6/XA9/MN1/a_324_334# 0.09fF
C2471 EN XA2/XA1/XA1/MP0/a_216_n18# 0.06fF
C2472 XA0/XA3/MP3/a_216_n18# D<8> 0.15fF
C2473 XDAC1/XC32a<0>/XRES2/B AVSS 3.96fF
C2474 XA0/XA3/MP2/a_216_n18# D<8> 0.15fF
C2475 XA7/XA5/MP3/a_216_n18# XA7/CN0 0.02fF
C2476 XA5/XA1/XA1/MP3/S XA20/CPO 0.01fF
C2477 XA5/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C2478 XA3/XA2/MP1/a_216_n18# XA3/XA2/MP2/a_216_n18# 0.01fF
C2479 XA0/XA6/MP0/a_216_n18# XA0/CN0 0.08fF
C2480 XA6/EN XA5/XA1/XA4/MN1/S 0.01fF
C2481 XA7/XA4/MN0/a_324_n18# AVSS 0.01fF
C2482 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC32a<0>/XRES16/B 0.05fF
C2483 XA8/XA11/A DONE 0.02fF
C2484 XDAC1/XC0/XRES8/B AVSS 9.01fF
C2485 XA20/CPO AVSS 5.39fF
C2486 XA20/XA2/MP0/a_216_n18# XA20/XA2/MP1/a_216_n18# 0.01fF
C2487 XDAC2/X16ab/XRES8/B AVSS 9.08fF
C2488 XA6/XA1/XA1/MP2/S XA6/XA1/XA1/MP3/G 0.04fF
C2489 XA5/XA1/XA4/MP1/a_216_n18# XA5/XA1/XA4/MP0/a_216_n18# 0.01fF
C2490 XA4/XA4/MN2/a_324_n18# XA4/XA4/MN1/a_324_n18# 0.01fF
C2491 XA1/XA2/MP0/a_216_n18# XA1/XA1/XA5/MP2/a_216_n18# 0.01fF
C2492 XA2/XA9/MN1/S XA2/XA9/Y 0.12fF
C2493 XA8/EN XA8/XA1/XA4/MN1/S 0.02fF
C2494 XA1/XA1/XA1/MP3/G XA20/CNO 0.06fF
C2495 XA6/XA9/B XA6/XA9/MN0/a_324_n18# 0.01fF
C2496 XA5/XA4/A VREF 0.37fF
C2497 XA2/XA1/XA4/MP2/a_216_n18# XA2/XA1/XA4/MP1/a_216_n18# 0.01fF
C2498 XA8/XA4/A XA20/XA3a/A 0.03fF
C2499 XA6/XA1/XA4/MN0/a_324_n18# XA6/XA1/XA4/MN1/a_324_n18# 0.01fF
C2500 XA1/XA2/MP1/a_216_n18# AVDD 0.08fF
C2501 XA20/XA3/N1 AVSS 0.93fF
C2502 D<7> VREF 1.73fF
C2503 XA3/XA1/XA5/MN2/S XA3/XA4/A 0.02fF
C2504 XA5/XA5/MN1/a_324_n18# XA5/XA5/MN2/a_324_n18# 0.01fF
C2505 VREF XA8/XA9/B 0.12fF
C2506 XA2/XA1/XA4/MP0/a_216_n18# XA2/XA1/XA2/MP0/a_216_n18# 0.01fF
C2507 XB1/XA5/MN1/a_324_334# AVSS 0.10fF
C2508 XA20/XA2/MP2/a_216_n18# AVDD 0.16fF
C2509 SARN XA20/XA3/CO 0.11fF
C2510 XA8/XA1/XA4/MN2/S AVSS 0.06fF
C2511 XA0/XA13/MP1/a_216_334# AVDD 0.17fF
C2512 XA3/CP0 XA3/XA5/MP0/a_216_n18# 0.07fF
C2513 D<3> XA5/XA3/MP1/a_216_n18# 0.03fF
C2514 XA2/EN XA1/XA9/A 0.09fF
C2515 XA0/XA1/XA1/MP3/G XA0/CN0 0.01fF
C2516 XDAC1/XC1/XRES1A/B XB1/XA4/GNG 0.76fF
C2517 VREF XA8/XA6/MP3/S 0.02fF
C2518 XA4/XA6/MP1/a_216_n18# D<4> 0.01fF
C2519 XA7/XA4/A XA7/CP0 0.52fF
C2520 XA7/XA3/MN0/a_324_n18# XA7/XA3/MN1/a_324_n18# 0.01fF
C2521 XA2/XA2/A XA2/XA1/XA5/MN2/S 0.05fF
C2522 XA5/XA5/MP2/a_216_n18# VREF 0.03fF
C2523 XA0/XA6/MP0/a_216_n18# XA0/XA5/MP3/a_216_n18# 0.01fF
C2524 XA4/XA4/MP1/a_216_n18# VREF 0.02fF
C2525 XA5/XA1/XA1/MN2/S AVDD 0.05fF
C2526 XB1/XA4/MN1/a_324_334# XB1/XA7/MN1/a_324_n18# 0.01fF
C2527 XA2/XA2/A XA2/XA2/MP0/a_216_n18# 0.08fF
C2528 XA4/XA1/XA5/MP2/a_216_n18# XA4/XA2/MP0/a_216_n18# 0.01fF
C2529 XA5/CP0 XA5/XA4/MN3/a_324_n18# 0.02fF
C2530 XDAC1/XC128a<1>/XRES16/B SARP 21.64fF
C2531 XA7/XA9/MP0/a_216_n18# AVDD 0.09fF
C2532 XA6/CN0 XA6/XA6/MP0/a_216_n18# 0.08fF
C2533 XA7/XA1/XA2/Y XA7/XA1/XA4/MN2/a_324_n18# 0.08fF
C2534 XA1/XA12/MP0/a_216_n18# XA1/XA12/A 0.07fF
C2535 XA2/XA4/MP2/a_216_n18# XA2/XA4/MP3/a_216_n18# 0.01fF
C2536 XA4/XA2/A XA4/XA2/MP2/a_216_n18# 0.15fF
C2537 XA4/XA2/MP0/a_216_n18# XA4/XA2/MP1/a_216_n18# 0.01fF
C2538 XB2/XA5/MP1/a_216_n18# XB2/XA5/MP1/a_216_334# 0.01fF
C2539 XA3/XA3/MN2/a_324_n18# XA3/CN1 0.16fF
C2540 D<8> XA0/CN0 2.94fF
C2541 XA7/XA9/Y AVSS 0.22fF
C2542 AVDD XA2/XA1/XA2/MP0/a_216_n18# 0.08fF
C2543 AVDD XA20/XA4/MP0/a_216_n18# 0.09fF
C2544 XA20/XA3/MN1/a_324_n18# XA20/XA3/N1 0.02fF
C2545 XA20/CPO XA0/XA1/XA1/MN2/a_324_n18# 0.08fF
C2546 XB2/XA3/B XA0/CEIN 0.01fF
C2547 XDAC2/XC128b<2>/XRES2/B SARN 3.05fF
C2548 D<4> XA1/CN0 0.05fF
C2549 XA4/XA9/Y AVDD 0.58fF
C2550 D<5> XA3/CP0 7.36fF
C2551 XA20/XA12/Y XA20/XA11/MP0/a_216_n18# 0.09fF
C2552 XA1/CP0 XA1/XA4/MN2/a_324_n18# 0.01fF
C2553 XA4/XA1/XA1/MP3/S AVDD 0.14fF
C2554 XA1/XA11/MP1/S AVDD 0.18fF
C2555 XA8/ENO XA20/CNO 0.27fF
C2556 XA6/CN1 XA6/XA3/MP1/a_216_n18# 0.15fF
C2557 XA4/XA1/XA1/MP3/G D<4> 0.02fF
C2558 XA6/XA5/MP2/a_216_n18# XA6/XA5/MP3/a_216_n18# 0.01fF
C2559 XA0/CEIN AVSS 3.81fF
C2560 XA1/XA9/A XA1/XA9/MN0/a_324_n18# 0.15fF
C2561 XA3/XA3/MP1/a_216_n18# VREF 0.02fF
C2562 XB1/XA0/MP0/a_216_n18# XB1/XA5b/MP1/a_216_n18# 0.01fF
C2563 EN XA0/XA2/MN0/a_324_n18# 0.07fF
C2564 XB2/M5/a_324_n18# XA0/CEIN 0.08fF
C2565 XA6/EN XA5/XA1/XA4/MP1/S 0.02fF
C2566 XB2/XA4/MN1/a_324_334# XB2/XA4/MN1/a_324_n18# 0.01fF
C2567 XA6/XA1/XA1/MP2/a_216_n18# XA6/XA1/XA1/MP1/a_216_n18# 0.01fF
C2568 XB2/M7/a_324_n18# SARP 0.02fF
C2569 XA6/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C2570 XA2/XA6/MP3/S AVDD 0.16fF
C2571 XA4/XA3/MP3/a_216_n18# D<4> 0.02fF
C2572 XB2/XA4/GNG XDAC2/XC1/XRES8/B 0.32fF
C2573 EN XA20/CPO 0.97fF
C2574 XA1/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C2575 XDAC1/XC0/XRES1B/B XDAC1/XC0/XRES4/B 1.64fF
C2576 XDAC1/XC0/XRES2/B XDAC1/XC0/XRES8/B 1.58fF
C2577 XA2/XA11/A XA2/CEO 0.02fF
C2578 XA3/XA2/MP0/a_216_n18# XA3/XA2/A 0.08fF
C2579 XDAC1/XC1/XRES8/B XDAC1/XC64a<0>/XRES16/B 0.03fF
C2580 XA8/ENO XA8/XA8/MP0/a_216_n18# 0.08fF
C2581 XA7/XA11/MN0/a_324_n18# XA7/XA9/Y 0.07fF
C2582 XDAC1/XC128b<2>/XRES16/B XDAC1/X16ab/XRES16/B 0.41fF
C2583 XA3/XA11/MP0/a_216_n18# XA3/XA11/MP1/a_216_n18# 0.01fF
C2584 XA6/EN XA5/XA2/A 0.10fF
C2585 AVDD XA0/XA1/XA1/MP2/S 0.11fF
C2586 XA2/CP0 XA1/CN0 0.05fF
C2587 XA4/XA9/Y XA4/XA9/MN1/S 0.12fF
C2588 XA5/XA1/XA4/MN0/a_324_n18# XA5/XA1/XA2/Y 0.02fF
C2589 XA4/CP0 XA3/CP0 0.03fF
C2590 XB2/CKN XB2/XA4/MN1/a_324_n18# 0.07fF
C2591 XB2/XA7/MN1/a_324_334# XB2/XA7/MN1/a_324_n18# 0.01fF
C2592 XA4/XA1/XA1/MN2/a_324_n18# XA4/XA1/XA1/MN1/a_324_n18# 0.01fF
C2593 XA5/XA1/XA4/MP2/a_216_n18# XA5/XA1/XA5/MP0/a_216_n18# 0.01fF
C2594 XA6/XA1/XA5/MN1/S XA20/CNO 0.01fF
C2595 XA5/XA1/XA2/MN0/a_324_n18# XA20/CPO 0.02fF
C2596 AVDD XA2/XA1/XA1/MP3/G 0.63fF
C2597 XA3/XA1/XA5/MP2/S XA4/EN 0.02fF
C2598 XA1/XA12/MP0/a_216_n18# XA1/XA13/MP1/a_216_n18# 0.01fF
C2599 XA2/XA1/XA4/MP2/S XA2/XA1/XA4/MN2/S 0.01fF
C2600 XA1/XA2/A XA0/XA2/A 0.03fF
C2601 XA20/XA2/MN5/a_324_n18# XA20/XA2/MN4/a_324_n18# 0.01fF
C2602 XA7/XA1/XA4/MN2/S XA7/EN 0.02fF
C2603 XA20/CNO XA2/XA1/XA1/MN2/a_324_n18# 0.07fF
C2604 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128a<1>/XRES2/B 1.58fF
C2605 XA0/XA5/MN0/a_324_n18# XA0/XA5/MN1/a_324_n18# 0.01fF
C2606 XA0/XA1/XA5/MN1/S AVSS 0.12fF
C2607 XA3/XA7/MP0/a_216_n18# XA4/EN 0.07fF
C2608 XA7/CEO XA8/XA9/Y 0.01fF
C2609 XDAC2/XC1/XRES8/B XDAC2/XC64a<0>/XRES1A/B 0.03fF
C2610 XA6/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C2611 XA2/EN XA1/XA2/A 0.10fF
C2612 EN XA0/XA1/XA5/MP1/S 0.04fF
C2613 XA4/XA6/MP0/a_216_n18# AVDD 0.08fF
C2614 XA4/XA1/XA1/MP2/a_216_n18# XA20/CNO 0.08fF
C2615 XA2/XA2/A XA4/EN 0.03fF
C2616 XA20/XA3a/A XA20/XA2a/MP1/a_216_n18# 0.01fF
C2617 XB1/XCAPB1/XCAPB4/m3_9756_132# XB1/XA3/B 0.07fF
C2618 XA2/XA1/XA1/MP3/S AVSS 0.02fF
C2619 AVDD XA2/XA13/MP1/a_216_n18# 0.13fF
C2620 XA7/XA8/MN0/a_324_n18# XA7/XA9/MN0/a_324_n18# 0.01fF
C2621 XA0/CP1 XA0/XA3/MP3/a_216_n18# 0.02fF
C2622 XA1/CP0 AVSS 1.73fF
C2623 XA20/XA11/MP0/a_216_n18# CK_SAMPLE 0.07fF
C2624 XA20/XA9/Y XA20/XA3/CO 0.34fF
C2625 XA0/CP1 XA0/XA3/MP2/a_216_n18# 0.01fF
C2626 XA4/XA9/MP1/a_216_n18# AVDD 0.09fF
C2627 XDAC2/XC64b<1>/XRES8/B XDAC2/X16ab/XRES8/B 0.21fF
C2628 XA3/XA1/XA5/MP1/S XA4/EN 0.02fF
C2629 XDAC2/X16ab/XRES1A/B XDAC2/X16ab/XRES16/B 1.60fF
C2630 EN XA5/XA1/XA4/MP0/a_216_n18# 0.07fF
C2631 XB2/XA7/MN1/a_324_334# XB2/XA2/MP0/G 0.07fF
C2632 D<4> XA4/XA3/MN3/a_324_n18# 0.02fF
C2633 XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C2634 XA0/XA5/MP0/a_216_n18# XA0/XA4/MP3/a_216_n18# 0.01fF
C2635 XA1/XA2/A XA1/XA2/MN0/a_324_n18# 0.08fF
C2636 XA20/XA4/MN1/a_324_n18# XA20/XA4/MP0/S 0.01fF
C2637 XA5/XA3/MP1/a_216_n18# XA5/XA3/MP2/a_216_n18# 0.01fF
C2638 XA1/XA4/A XA20/CNO 0.21fF
C2639 XA2/CP0 XA3/EN 0.12fF
C2640 XB2/M8/a_324_334# SARP 0.01fF
C2641 XA7/XA4/MP3/a_216_n18# AVDD 0.07fF
C2642 XDAC2/XC64b<1>/XRES1A/B XDAC2/X16ab/XRES1B/B 0.63fF
C2643 XA2/CEO AVSS 0.46fF
C2644 XDAC2/XC128a<1>/XRES2/B SARN 3.05fF
C2645 XA6/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C2646 XB1/XA4/GNG XB1/XA4/MN1/S 0.01fF
C2647 XA8/XA3/MN3/a_324_n18# XA8/XA4/A 0.01fF
C2648 XA2/CN0 XA2/XA2/A 0.03fF
C2649 XA7/XA1/XA1/MP2/a_216_n18# XA20/CPO 0.06fF
C2650 XA1/XA1/XA5/MN2/a_324_n18# XA1/XA1/XA2/Y 0.07fF
C2651 XB1/XA5/MN1/a_324_n18# XB1/XA5/MN1/a_324_334# 0.01fF
C2652 XA20/CNO XA20/XA3a/MP1/a_216_n18# 0.01fF
C2653 XA5/XA1/XA1/MN2/S XA5/EN 0.05fF
C2654 CK_SAMPLE_BSSW XB1/XA4/GNG 0.03fF
C2655 EN XA0/XA1/XA5/MP0/a_216_n18# 0.16fF
C2656 XA4/XA5/MN2/a_324_n18# XA4/XA5/MN3/a_324_n18# 0.01fF
C2657 XA7/XA12/MP0/a_216_n18# XA6/CEO 0.08fF
C2658 XB1/XCAPB1/XCAPB2/m3_252_308# XB1/XA3/B 0.02fF
C2659 D<6> D<8> 0.07fF
C2660 XA4/XA1/XA5/MP1/S AVDD 0.13fF
C2661 XA7/XA1/XA2/Y XA7/XA1/XA5/MN1/S 0.05fF
C2662 XA0/XA4/A D<8> 0.62fF
C2663 XA0/CP0 XA20/CNO 0.05fF
C2664 XA7/XA3/MP2/a_216_n18# XA7/CN1 0.15fF
C2665 XA6/XA4/MP1/a_216_n18# XA6/XA4/MP2/a_216_n18# 0.01fF
C2666 XA20/XA9/A XA20/XA3/CO 0.22fF
C2667 AVDD XA3/XA4/A 1.42fF
C2668 XA7/XA1/XA5/MN2/a_324_n18# XA7/XA2/MN0/a_324_n18# 0.01fF
C2669 EN XA0/XA1/XA4/MN2/a_324_n18# 0.08fF
C2670 XA4/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C2671 XA8/XA9/A XA8/XA9/B 0.29fF
C2672 XA0/CEO AVDD 1.51fF
C2673 XA0/XA1/XA4/MN2/S XA0/XA1/XA4/MN1/S 0.04fF
C2674 XA5/CN1 XA4/CN1 0.03fF
C2675 XA2/XA4/A D<6> 0.26fF
C2676 XDAC2/XC64b<1>/XRES4/B XDAC2/XC64b<1>/XRES16/B 0.25fF
C2677 XA6/EN XA5/XA1/XA5/MP1/S 0.02fF
C2678 XA6/CN0 AVDD 5.33fF
C2679 XA0/XA3/MP0/a_216_n18# VREF 0.02fF
C2680 XA4/XA1/XA1/MP3/S XA5/EN 0.10fF
C2681 XA2/XA9/MP0/a_216_n18# XA2/XA9/A 0.14fF
C2682 XDAC1/XC1/XRES4/B XDAC1/XC1/XRES2/B 0.55fF
C2683 XA7/XA9/B XA7/XA9/A 0.29fF
C2684 XA1/XA1/XA5/MP0/a_216_n18# XA1/XA1/XA4/MP2/a_216_n18# 0.01fF
C2685 XA1/XA4/MP3/a_216_n18# AVDD 0.07fF
C2686 XA5/XA11/MN1/a_324_n18# AVSS 0.01fF
C2687 XA20/XA4/MN1/a_324_n18# XA20/XA4/MN0/a_324_n18# 0.01fF
C2688 XA1/XA2/MP3/a_216_n18# VREF 0.03fF
C2689 XA3/XA9/A XA3/XA9/B 0.29fF
C2690 XA3/XA1/XA1/MP2/S XA3/XA1/XA1/MP3/G 0.04fF
C2691 XA5/XA13/MP1/a_216_334# XA5/XA13/MP1/a_216_n18# 0.01fF
C2692 XA6/EN XA5/CN1 0.10fF
C2693 XA4/XA11/A XA4/XA11/MP0/a_216_n18# 0.07fF
C2694 XA7/XA1/XA2/Y XA7/XA1/XA4/MN0/a_324_n18# 0.02fF
C2695 XA20/CNO XA0/XA1/XA1/MN1/a_324_n18# 0.07fF
C2696 XA8/XA11/MN0/a_324_n18# XA8/XA9/Y 0.07fF
C2697 XA0/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C2698 XA8/EN XA8/XA4/A 0.14fF
C2699 XA6/XA1/XA2/Y AVDD 0.33fF
C2700 XA1/CP0 CK_SAMPLE 0.09fF
C2701 XDAC2/XC1/XRES16/B SARN 21.64fF
C2702 XA20/XA3/N2 VREF 0.01fF
C2703 XA20/XA3/MN5/a_324_n18# XA20/XA3/MN4/a_324_n18# 0.01fF
C2704 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128b<2>/XRES4/B 0.29fF
C2705 XDAC2/XC128b<2>/XRES2/B XDAC2/XC128b<2>/XRES1B/B 0.23fF
C2706 AVDD XB1/XA5/MP1/a_216_334# 0.17fF
C2707 XA3/XA2/A VREF 0.36fF
C2708 EN XA0/XA1/XA5/MN1/S 0.02fF
C2709 XB1/XCAPB1/XCAPB3/m3_9756_132# XB1/XA4/GNG 0.02fF
C2710 XA5/XA6/MN2/a_324_n18# AVSS 0.01fF
C2711 XA0/CP1 XA0/CN0 0.46fF
C2712 D<8> SARP 0.09fF
C2713 XA7/XA1/XA5/MP0/a_216_n18# XA7/XA1/XA5/MP1/a_216_n18# 0.01fF
C2714 XA8/XA7/MP0/a_216_n18# XA8/XA6/MP3/a_216_n18# 0.01fF
C2715 VREF XA8/CP0 0.71fF
C2716 D<3> XA5/XA6/MP3/S 0.02fF
C2717 XA20/XA11/MP1/S XA20/XA11/Y 0.07fF
C2718 XA1/CP0 EN 0.05fF
C2719 XA6/XA7/MN0/a_324_n18# XA6/XA6/MN3/a_324_n18# 0.01fF
C2720 XDAC2/XC1/XRES1B/B XDAC2/XC1/XRES16/B 0.12fF
C2721 XDAC2/XC0/XRES8/B AVSS 9.01fF
C2722 XA3/XA4/MP0/a_216_n18# VREF 0.02fF
C2723 XDAC2/XC128a<1>/XRES1A/B XDAC2/XC32a<0>/XRES16/B 0.04fF
C2724 XA0/XA12/A XA0/XA12/MP0/a_216_n18# 0.07fF
C2725 XA7/XA4/MP2/a_216_n18# AVDD 0.07fF
C2726 XA6/CP0 XA6/XA4/MP1/a_216_n18# 0.02fF
C2727 XA7/XA1/XA2/Y XA20/CNO 0.22fF
C2728 XA1/XA2/MP1/a_216_n18# XA1/XA2/A 0.15fF
C2729 XA6/XA1/XA4/MN1/S XA6/XA4/A 0.02fF
C2730 XA6/XA6/MN0/a_324_n18# XA6/XA6/MN1/a_324_n18# 0.01fF
C2731 XA4/XA4/A XA20/CNO 0.18fF
C2732 XA0/XA1/XA5/MP2/S AVDD 0.08fF
C2733 VREF XA8/XA9/A 0.03fF
C2734 XA5/XA9/Y XA5/XA12/A 0.02fF
C2735 XA1/XA1/XA5/MN1/S XA20/CNO 0.01fF
C2736 XA5/XA4/MN0/a_324_n18# XA5/XA4/MN1/a_324_n18# 0.01fF
C2737 XB2/XA7/MP1/a_216_n18# AVDD 0.15fF
C2738 XA8/XA6/MN0/a_324_n18# AVSS 0.01fF
C2739 XA6/XA5/MN0/a_324_n18# XA6/XA4/A 0.07fF
C2740 XA2/EN XA1/CN1 0.25fF
C2741 XA1/XA6/MP0/a_216_n18# AVDD 0.08fF
C2742 XA4/EN XA3/XA1/XA2/Y 0.14fF
C2743 XA4/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C2744 XA6/XA2/A XA20/CNO 0.03fF
C2745 XA20/CPO XA6/XA1/XA1/MP3/G 0.14fF
C2746 XA5/XA9/MN1/a_324_334# XA5/XA11/MN0/a_324_n18# 0.01fF
C2747 XA0/XA2/MN2/a_324_n18# D<8> 0.02fF
C2748 XA2/XA1/XA2/Y XA2/XA1/XA4/MP1/S 0.01fF
C2749 D<0> XA8/XA4/A 0.22fF
C2750 XA6/XA1/XA1/MP2/a_216_n18# XA6/XA1/XA1/MP3/G 0.01fF
C2751 XA2/XA12/A XA2/CEO 0.11fF
C2752 XA7/XA1/XA1/MP3/S XA7/XA1/XA1/MP3/G 0.04fF
C2753 XA6/XA1/XA5/MP2/S EN 0.04fF
C2754 XA3/CP0 AVDD 1.48fF
C2755 XA20/XA3/N1 XA20/XA3/MN3/a_324_n18# 0.02fF
C2756 XA5/XA12/A XA5/XA11/A 0.07fF
C2757 XA20/XA12/MP0/a_216_n18# DONE 0.08fF
C2758 XA4/XA2/A VREF 0.36fF
C2759 XA20/XA3/MP6/a_216_n18# XA20/XA3a/A 0.15fF
C2760 XDAC2/XC128b<2>/XRES16/B SARN 21.64fF
C2761 XA2/XA4/A XA2/XA4/MN0/a_324_n18# 0.09fF
C2762 XDAC2/XC64b<1>/XRES4/B SARN 6.32fF
C2763 AVSS XA8/XA9/Y 0.22fF
C2764 XA5/XA2/MN2/a_324_n18# AVSS 0.01fF
C2765 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MP2/a_216_n18# 0.01fF
C2766 XA5/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C2767 XA4/XA1/XA5/MP1/S XA5/EN 0.02fF
C2768 XA7/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C2769 VREF XA2/XA4/MP2/a_216_n18# 0.03fF
C2770 XA7/XA9/A AVSS 0.31fF
C2771 XDAC1/XC128b<2>/XRES1B/B XDAC1/X16ab/XRES16/B 0.05fF
C2772 XA3/CN0 XA3/XA6/MP2/a_216_n18# 0.08fF
C2773 XDAC2/XC64a<0>/XRES1A/B XDAC2/XC64a<0>/XRES16/B 1.60fF
C2774 XA5/XA1/XA1/MN1/a_324_n18# XA5/XA1/XA1/MN2/a_324_n18# 0.01fF
C2775 XB2/CKN XB2/M4/G 0.28fF
C2776 XB2/XA7/MN1/a_324_n18# XB2/XA1/MP0/G 0.07fF
C2777 D<7> XA1/XA3/MP2/a_216_n18# 0.01fF
C2778 XDAC2/XC128b<2>/XRES4/B XDAC2/XC128a<1>/XRES4/B 0.10fF
C2779 XA8/XA12/A XA8/XA13/MN1/a_324_n18# 0.07fF
C2780 XDAC2/XC128a<1>/XRES16/B SARN 21.64fF
C2781 XA2/EN XA1/XA8/MP0/a_216_n18# 0.08fF
C2782 XA0/XA4/A XA0/XA1/XA5/MN2/S 0.02fF
C2783 XA0/XA6/MN1/S AVSS 0.15fF
C2784 XA1/XA1/XA5/MP0/a_216_n18# EN 0.16fF
C2785 XA4/XA1/XA4/MP1/S EN 0.02fF
C2786 SAR_IP XA0/CEIN 0.33fF
C2787 XA7/CP0 XA7/EN 0.03fF
C2788 XA20/XA3/N2 XA20/XA4/MP0/S 0.01fF
C2789 XA5/XA1/XA1/MN1/a_324_n18# AVSS 0.01fF
C2790 AVDD XA3/XA4/MP1/a_216_n18# 0.07fF
C2791 XA7/XA6/MN1/a_324_n18# XA7/XA6/MN0/a_324_n18# 0.01fF
C2792 XA2/CN1 XA20/CPO 0.18fF
C2793 XA1/XA11/MN1/a_324_n18# XA0/CEO 0.08fF
C2794 D<7> XDAC1/XC64b<1>/XRES16/B 0.17fF
C2795 XA8/XA3/MN2/a_324_n18# XA8/XA4/A 0.01fF
C2796 XA6/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C2797 EN XA0/XA1/XA4/MP2/S 0.03fF
C2798 XA8/XA1/XA1/MP1/a_216_n18# AVDD 0.08fF
C2799 XB1/XCAPB1/XCAPB3/m3_9828_132# XB1/XA3/B 0.21fF
C2800 XA8/XA2/MN1/a_324_n18# XA8/XA2/A 0.15fF
C2801 XA4/XA3/MP1/a_216_n18# XA4/CN1 0.15fF
C2802 XA4/XA1/XA5/MP2/S AVDD 0.08fF
C2803 CK_SAMPLE XA8/XA6/MN0/a_324_n18# 0.08fF
C2804 XA6/XA1/XA2/Y XA5/EN 0.02fF
C2805 XA0/CP1 D<6> 1.34fF
C2806 D<2> XA6/XA1/XA1/MN2/S 0.02fF
C2807 XB2/XA2/MP0/G XB2/XA1/MP0/G 0.02fF
C2808 XA0/CP1 XA0/XA4/A 0.26fF
C2809 XA7/XA4/MP1/a_216_n18# AVDD 0.07fF
C2810 XA1/XA4/A XA1/XA3/MN2/a_324_n18# 0.01fF
C2811 D<2> XA6/XA3/MN1/a_324_n18# 0.02fF
C2812 XA2/CN0 XA2/XA5/MN1/a_324_n18# 0.02fF
C2813 XA2/XA9/MP1/a_216_n18# AVDD 0.09fF
C2814 XDAC2/XC64b<1>/XRES16/B XA0/CN0 0.02fF
C2815 XA3/XA1/XA4/MN2/S XA4/EN 0.01fF
C2816 XA7/XA1/XA1/MP3/G AVSS 0.12fF
C2817 XA2/XA4/A XA2/XA4/MN1/a_324_n18# 0.15fF
C2818 XA8/XA1/XA2/Y XA8/XA1/XA5/MN2/a_324_n18# 0.07fF
C2819 XA1/XA3/MP1/a_216_n18# D<7> 0.02fF
C2820 XA3/XA5/MN1/a_324_n18# XA3/XA5/MN0/a_324_n18# 0.01fF
C2821 XA6/EN XA7/EN 0.06fF
C2822 XA3/CN0 XA3/XA6/MP0/a_216_n18# 0.08fF
C2823 XA5/XA1/XA1/MP3/G XA20/CPO 0.15fF
C2824 XA6/XA1/XA2/MN0/a_324_n18# XA6/XA1/XA1/MP3/G 0.06fF
C2825 XA8/XA3/MN1/a_324_n18# XA8/XA3/MN0/a_324_n18# 0.01fF
C2826 XA8/XA13/MP1/a_216_334# XA8/XA13/MP1/a_216_n18# 0.01fF
C2827 XB2/XA2/MP0/G XB2/XA7/MP1/a_216_334# 0.07fF
C2828 XA2/EN XA1/XA7/MN0/a_324_n18# 0.08fF
C2829 CK_SAMPLE XA8/XA9/Y 0.01fF
C2830 XA6/XA9/A XA6/XA8/MP0/a_216_n18# 0.07fF
C2831 XA5/XA3/MN3/a_324_n18# XA5/CN1 0.15fF
C2832 XDAC2/XC64a<0>/XRES1B/B AVSS 3.58fF
C2833 XDAC2/X16ab/XRES16/B D<8> 0.05fF
C2834 XA8/XA3/MP2/a_216_n18# XA8/XA3/MP3/a_216_n18# 0.01fF
C2835 XA6/XA6/MN3/S AVSS 0.13fF
C2836 XA2/XA1/XA5/MN1/S AVSS 0.12fF
C2837 D<5> XA3/XA7/MP0/a_216_n18# 0.08fF
C2838 XA7/XA9/A CK_SAMPLE 0.02fF
C2839 XA7/XA1/XA5/MP2/a_216_n18# EN 0.16fF
C2840 XA5/XA12/A XA5/CEO 0.20fF
C2841 XA1/XA3/MP2/a_216_n18# VREF 0.03fF
C2842 EN XA2/XA1/XA5/MP1/S 0.03fF
C2843 XA7/XA5/MP2/a_216_n18# AVDD 0.07fF
C2844 XA0/XA6/MN1/S CK_SAMPLE 0.04fF
C2845 XA5/XA5/MP1/a_216_n18# XA5/CN0 0.02fF
C2846 XA1/XA2/MP1/a_216_n18# XA1/CN1 0.02fF
C2847 XA4/CN0 D<8> 0.07fF
C2848 XA3/XA3/MN0/a_324_n18# XA3/XA2/A 0.07fF
C2849 XDAC2/XC0/XRES1A/B XDAC2/XC0/XRES8/B 0.12fF
C2850 XA20/XA3/MP1/a_216_n18# XA20/XA3/MP0/a_216_n18# 0.01fF
C2851 XA0/XA12/A AVSS 0.41fF
C2852 XDAC2/XC64b<1>/XRES8/B XDAC2/XC0/XRES8/B 0.21fF
C2853 XA7/XA3/MP1/a_216_n18# XA7/XA3/MP0/a_216_n18# 0.01fF
C2854 XA5/CEO XA6/XA11/MP1/a_216_n18# 0.06fF
C2855 XDAC2/XC128b<2>/XRES8/B XDAC2/X16ab/XRES8/B 0.21fF
C2856 XA7/XA9/MP1/a_216_334# XA7/XA11/MP0/a_216_n18# 0.01fF
C2857 XDAC2/XC64a<0>/XRES2/B XDAC2/XC64a<0>/XRES4/B 0.55fF
C2858 XA0/CP1 SARP 0.61fF
C2859 XA0/XA1/XA4/MN1/S XA0/XA1/XA4/MP1/S 0.01fF
C2860 XA5/XA4/A XA20/CPO 0.03fF
C2861 XDAC2/XC32a<0>/XRES1B/B XDAC2/XC32a<0>/XRES8/B 0.12fF
C2862 XB2/XA1/Y XB2/XA3/B 0.01fF
C2863 XA5/XA1/XA1/MP2/S AVDD 0.09fF
C2864 D<7> XA20/CPO 0.06fF
C2865 XA8/XA9/MN0/a_324_n18# XA8/XA9/B 0.01fF
C2866 XA5/CN0 D<8> 0.06fF
C2867 XA7/CN1 XA8/XA4/A 0.04fF
C2868 XA6/CN0 XDAC2/XC32a<0>/XRES16/B 0.02fF
C2869 XB2/XA1/Y AVSS 0.33fF
C2870 XA8/ENO XA8/XA4/A 0.11fF
C2871 XA20/CNO XA2/XA1/XA5/MN1/a_324_n18# 0.07fF
C2872 XA5/XA11/MP1/S XA4/CEO 0.02fF
C2873 XB2/XCAPB1/XCAPB4/m3_252_308# XB2/XA4/GNG 0.13fF
C2874 XA5/XA13/MN1/a_324_n18# AVSS 0.09fF
C2875 XA20/XA3a/MN2/a_324_n18# XA20/XA3a/MN3/a_324_n18# 0.01fF
C2876 XA8/XA2/MN3/a_324_n18# XA8/XA2/A 0.15fF
C2877 XB2/M4/G XA0/CEIN 0.27fF
C2878 XA3/XA2/MP3/a_216_n18# XA3/XA3/MP0/a_216_n18# 0.01fF
C2879 XDAC2/XC1/XRES4/B XDAC2/XC1/XRES8/B 2.60fF
C2880 XB2/XA4/MN1/a_324_334# XB2/XA1/MP0/G 0.08fF
C2881 XA0/XA9/MN1/S AVDD 0.01fF
C2882 D<7> XA1/XA7/MP0/a_216_n18# 0.08fF
C2883 XA3/XA1/XA5/MP2/S XA3/XA1/XA5/MN2/S 0.01fF
C2884 XDAC1/XC64a<0>/XRES8/B AVSS 9.11fF
C2885 XA0/XA4/A XA0/XA1/XA4/MN1/S 0.02fF
C2886 CK_SAMPLE_BSSW XB1/XA3/MP0/S 0.01fF
C2887 XA2/CN0 XA0/CN0 1.01fF
C2888 XA3/XA2/A XA4/XA2/A 0.03fF
C2889 XA6/XA9/MN1/S AVSS 0.15fF
C2890 XA5/XA1/XA1/MP3/a_216_n18# AVDD 0.08fF
C2891 AVDD XA20/XA3/CO 4.14fF
C2892 XA1/XA3/MP1/a_216_n18# VREF 0.02fF
C2893 XB2/XCAPB1/XCAPB0/m3_9756_132# XB2/XA3/B 0.07fF
C2894 XA20/XA3a/MN1/a_324_n18# XA20/XA3a/A 0.15fF
C2895 XA0/XA9/Y VREF 0.03fF
C2896 XA4/XA1/XA5/MP2/a_216_n18# EN 0.16fF
C2897 XA5/XA12/MN0/a_324_n18# XA4/CEO 0.07fF
C2898 XA5/XA1/XA5/MN1/S AVDD 0.02fF
C2899 XA3/XA13/MP1/a_216_n18# XA3/XA12/MP0/a_216_n18# 0.01fF
C2900 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC64b<1>/XRES8/B 0.12fF
C2901 XA0/XA9/A XA1/EN 0.09fF
C2902 XA3/EN XA2/XA1/XA1/MN2/S 0.06fF
C2903 XA4/XA1/XA5/MP1/S XA4/XA1/XA5/MN1/S 0.01fF
C2904 XDAC2/XC64b<1>/XRES16/B XDAC2/X16ab/XRES2/B 0.01fF
C2905 XA1/XA6/MP1/a_216_n18# AVDD 0.08fF
C2906 XA0/CP0 XA0/XA5/MN2/a_324_n18# 0.15fF
C2907 XA7/XA6/MN3/a_324_n18# XA7/XA7/MN0/a_324_n18# 0.01fF
C2908 XA7/XA1/XA4/MP0/a_216_n18# EN 0.07fF
C2909 D<1> D<4> 0.05fF
C2910 XA0/XA4/A XA0/XA3/MN3/a_324_n18# 0.01fF
C2911 XA8/CN0 XA8/XA5/MP1/a_216_n18# 0.02fF
C2912 XA3/XA1/XA5/MN1/S XA3/XA1/XA5/MN2/S 0.04fF
C2913 XA6/XA9/B AVSS 0.61fF
C2914 XA6/XA2/MP3/a_216_n18# VREF 0.03fF
C2915 XDAC2/XC128b<2>/XRES1B/B XDAC2/XC128b<2>/XRES16/B 0.12fF
C2916 XA20/XA2/MN6/a_324_334# XA20/XA2a/MN1/a_324_n18# 0.01fF
C2917 XDAC1/XC128a<1>/XRES2/B AVSS 3.71fF
C2918 XA0/XA9/MN1/a_324_n18# XA0/XA9/MN1/a_324_334# 0.01fF
C2919 XA6/XA1/XA5/MN2/S XA20/CNO 0.01fF
C2920 XA7/XA1/XA1/MP3/G EN 0.10fF
C2921 XB2/CKN XB2/XA1/MP0/G 0.03fF
C2922 XA3/XA1/XA4/MN1/a_324_n18# XA3/XA1/XA4/MN0/a_324_n18# 0.01fF
C2923 XA7/XA3/MN0/a_324_n18# XA7/XA2/A 0.07fF
C2924 XA6/XA6/MN3/S CK_SAMPLE 0.03fF
C2925 XA7/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C2926 SARN XA0/CN0 0.80fF
C2927 XA4/CN0 XA4/CN1 0.08fF
C2928 XA7/XA6/MP2/a_216_n18# XA7/XA6/MP3/a_216_n18# 0.01fF
C2929 AVDD XB1/XA2/MP0/G 0.45fF
C2930 XA7/XA1/XA0/MP1/a_216_n18# XA7/XA1/XA1/MP0/a_216_n18# 0.01fF
C2931 XA8/XA4/A XA8/CN0 0.03fF
C2932 XA0/XA4/MP0/a_216_n18# VREF 0.02fF
C2933 XA6/XA1/XA5/MN1/a_324_n18# XA6/XA1/XA5/MN0/a_324_n18# 0.01fF
C2934 XB2/XCAPB1/XCAPB2/m3_9756_132# XB2/XA4/GNG 0.02fF
C2935 XA20/XA2/MP4/a_216_n18# XA20/XA2/MP5/a_216_n18# 0.01fF
C2936 XA5/EN XA4/XA1/XA5/MP2/S 0.02fF
C2937 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC32a<0>/XRES8/B 0.12fF
C2938 XA8/ENO XA8/XA1/XA2/MN0/a_324_n18# 0.09fF
C2939 XA3/XA9/A AVSS 0.31fF
C2940 XA20/XA1/MP6_DMY/a_216_n18# AVDD 0.24fF
C2941 XA6/EN XA4/CN0 0.04fF
C2942 XA6/XA9/Y XA6/XA9/MN1/S 0.12fF
C2943 XA6/XA4/A XA7/XA4/A 0.03fF
C2944 XA6/XA9/B XA5/XA9/B 0.07fF
C2945 XA7/XA5/MN3/a_324_n18# XA7/XA6/MN0/a_324_n18# 0.01fF
C2946 EN XA2/XA1/XA5/MN1/S 0.01fF
C2947 VREF XA20/CPO 0.03fF
C2948 XA1/CP0 XA2/CN1 0.10fF
C2949 XA8/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C2950 XA5/XA3/MP3/a_216_n18# AVDD 0.07fF
C2951 XA2/XA8/MP0/a_216_n18# XA2/XA7/MP0/a_216_n18# 0.01fF
C2952 XA4/XA9/B XA4/XA6/MP3/S 0.07fF
C2953 XB1/M4/G XB1/M4/a_324_n18# 0.15fF
C2954 XA2/XA4/MN2/a_324_n18# AVSS 0.01fF
C2955 XA2/XA5/MP2/a_216_n18# XA2/XA5/MP1/a_216_n18# 0.01fF
C2956 XA0/XA2/A AVSS 0.22fF
C2957 XA4/CN1 XA4/XA4/MN0/a_324_n18# 0.07fF
C2958 XB2/M8/a_324_n18# SARP 0.02fF
C2959 XA4/XA1/XA4/MP2/S XA4/XA4/A 0.05fF
C2960 XA6/EN XA5/CN0 0.20fF
C2961 XA3/CEO XA4/CEO 0.03fF
C2962 XDAC1/XC32a<0>/XRES4/B XDAC1/XC128a<1>/XRES4/B 0.10fF
C2963 XA8/XA12/A AVDD 0.45fF
C2964 XA0/XA9/A XA0/DONE 0.07fF
C2965 XA2/EN XA1/XA6/MP3/S 0.02fF
C2966 XA2/XA5/MN1/a_324_n18# XA2/XA5/MN2/a_324_n18# 0.01fF
C2967 XA6/XA4/A XA5/XA2/A 0.03fF
C2968 XA2/EN AVSS 1.36fF
C2969 XA7/XA5/MN2/a_324_n18# XA7/CP0 0.15fF
C2970 XA6/XA9/B XA6/XA9/Y 0.15fF
C2971 XA6/XA3/MN0/a_324_n18# XA6/XA2/MN3/a_324_n18# 0.01fF
C2972 XA20/XA13/MP1/a_216_n18# XA20/XA12/MP0/a_216_n18# 0.01fF
C2973 XA1/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C2974 XA20/XA3/MP3/a_216_n18# XA20/XA9/Y 0.07fF
C2975 XA4/XA7/MP0/a_216_n18# D<4> 0.08fF
C2976 XA20/CNO XA0/XA1/XA2/Y 0.21fF
C2977 D<4> XA3/CN1 0.23fF
C2978 XA8/XA9/Y XA8/XA9/MN1/S 0.12fF
C2979 XA5/XA12/MP0/a_216_n18# AVDD 0.08fF
C2980 D<2> XA6/XA7/MP0/a_216_n18# 0.08fF
C2981 XA3/XA5/MN3/a_324_n18# XA3/CP0 0.15fF
C2982 XA5/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C2983 AVDD XA2/XA1/XA5/MP2/S 0.08fF
C2984 XA7/CN0 XA7/XA6/MP0/a_216_n18# 0.08fF
C2985 XA3/XA8/MN0/a_324_n18# XA3/XA9/MN0/a_324_n18# 0.01fF
C2986 XDAC1/XC128b<2>/XRES4/B XDAC1/X16ab/XRES16/B 0.03fF
C2987 XA1/XA1/XA1/MP1/a_216_n18# XA1/XA1/XA1/MP2/a_216_n18# 0.01fF
C2988 D<6> XA4/EN 0.02fF
C2989 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC0/XRES1A/B 0.63fF
C2990 XA4/XA3/MN2/a_324_n18# XA4/CN1 0.16fF
C2991 XA5/XA1/XA4/MN0/a_324_n18# XA5/XA1/XA4/MN1/a_324_n18# 0.01fF
C2992 D<5> XA3/XA1/XA2/Y 0.02fF
C2993 XA1/EN AVDD 4.88fF
C2994 XA7/XA6/MN1/S AVDD 0.01fF
C2995 XB1/XCAPB1/XCAPB0/m3_9756_132# XB1/XA4/GNG 0.02fF
C2996 XA6/XA9/B CK_SAMPLE 0.09fF
C2997 XA0/XA1/XA5/MP1/S VREF 0.02fF
C2998 XA8/EN XA8/XA1/XA1/MP3/G 0.03fF
C2999 XA5/XA1/XA1/MP2/S XA5/EN 0.01fF
C3000 D<2> D<4> 0.66fF
C3001 XA6/CP0 XA7/CP0 0.03fF
C3002 XA1/CEO XA2/XA11/MP1/a_216_n18# 0.06fF
C3003 XA2/XA2/A XA2/XA2/MP2/a_216_n18# 0.15fF
C3004 XA3/XA2/MP1/a_216_n18# AVDD 0.08fF
C3005 XA6/XA2/A XA6/XA2/MN2/a_324_n18# 0.15fF
C3006 XA7/XA1/XA1/MP2/a_216_n18# XA7/XA1/XA1/MP3/G 0.01fF
C3007 XA6/XA11/MP1/S XA6/XA12/A 0.06fF
C3008 XA8/XA1/XA2/Y XA20/CPO 0.22fF
C3009 XA0/XA1/XA1/MN3/a_324_n18# XA0/XA1/XA1/MN2/a_324_n18# 0.01fF
C3010 XA1/XA12/A XA1/CEO 0.20fF
C3011 XA8/EN XA7/XA1/XA5/MP2/S 0.02fF
C3012 XA3/XA1/XA4/MP1/S XA3/XA1/XA2/Y 0.01fF
C3013 XA1/CEO XA2/XA11/MN1/a_324_n18# 0.08fF
C3014 XA8/XA12/MN0/a_324_n18# XA8/XA13/MN1/a_324_n18# 0.01fF
C3015 XDAC2/XC64b<1>/XRES1A/B AVSS 2.95fF
C3016 XA1/XA3/MN3/a_324_n18# XA1/XA3/MN2/a_324_n18# 0.01fF
C3017 XA2/CP0 XA3/CN1 0.10fF
C3018 XA6/CN1 D<1> 0.01fF
C3019 XA2/CN0 D<6> 0.46fF
C3020 XDAC2/X16ab/XRES2/B SARN 3.05fF
C3021 XA7/XA9/Y VREF 0.03fF
C3022 XA3/XA1/XA4/MP2/S XA4/EN 0.02fF
C3023 XA3/XA9/A CK_SAMPLE 0.02fF
C3024 XA8/XA5/MP0/a_216_n18# XA8/XA5/MP1/a_216_n18# 0.01fF
C3025 XA8/XA6/MP2/a_216_n18# XA8/XA6/MP1/a_216_n18# 0.01fF
C3026 XA5/XA7/MP0/a_216_n18# XA6/EN 0.07fF
C3027 XDAC1/XC1/XRES2/B XDAC1/XC64a<0>/XRES16/B 0.01fF
C3028 XA4/XA9/MP0/a_216_n18# AVDD 0.09fF
C3029 XA20/XA1/MN2/a_324_n18# SARP 0.15fF
C3030 XA1/CP0 D<7> 5.63fF
C3031 D<3> D<4> 3.24fF
C3032 XB2/XA1/Y XB2/XA4/MN1/a_324_n18# 0.08fF
C3033 XA7/XA1/XA4/MP2/S XA7/XA1/XA4/MN2/S 0.01fF
C3034 XA20/XA10/MN1/S AVSS 0.12fF
C3035 XDAC2/XC128a<1>/XRES2/B XDAC2/XC32a<0>/XRES2/B 0.05fF
C3036 XA0/XA9/MN1/a_324_334# XA0/XA11/MN0/a_324_n18# 0.01fF
C3037 XA7/XA1/XA1/MN1/a_324_n18# XA7/XA1/XA1/MN2/a_324_n18# 0.01fF
C3038 VREF XA0/CEIN 0.05fF
C3039 XB2/XA1/MP0/G XA0/CEIN 0.04fF
C3040 XA2/XA1/XA2/Y XA2/XA1/XA5/MN1/a_324_n18# 0.09fF
C3041 XA8/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C3042 XA8/XA1/XA2/Y XA8/XA1/XA4/MN2/S 0.05fF
C3043 XDAC1/XC1/XRES8/B XDAC1/XC1/XRES1B/B 0.12fF
C3044 XA8/XA5/MP0/a_216_n18# XA8/XA4/A 0.08fF
C3045 XA1/XA1/XA1/MN2/S AVSS 0.27fF
C3046 XA1/XA1/XA1/MP2/S XA1/XA1/XA1/MP3/G 0.04fF
C3047 XA2/XA1/XA4/MP2/a_216_n18# XA2/XA1/XA5/MP0/a_216_n18# 0.01fF
C3048 XA2/EN CK_SAMPLE 0.09fF
C3049 D<6> SARN 0.03fF
C3050 XA6/CN0 XA1/CN1 0.05fF
C3051 XA0/DONE AVDD 0.21fF
C3052 XA0/XA2/A EN 0.22fF
C3053 XA2/XA4/MN3/a_324_n18# XA2/XA4/MN2/a_324_n18# 0.01fF
C3054 XA3/XA11/MP1/a_216_n18# XA3/XA12/MP0/a_216_n18# 0.01fF
C3055 XA5/XA1/XA1/MP3/a_216_n18# XA5/XA1/XA2/MP0/a_216_n18# 0.01fF
C3056 XA0/XA1/XA5/MN0/a_324_n18# XA0/XA1/XA4/MN2/a_324_n18# 0.01fF
C3057 XA3/XA5/MN0/a_324_n18# XA3/XA4/MN3/a_324_n18# 0.01fF
C3058 XA5/XA1/XA2/Y AVDD 0.33fF
C3059 XA8/XA4/MN2/a_324_n18# XA8/XA4/A 0.15fF
C3060 XA20/XA1/MP2_DMY/a_216_n18# AVDD 0.24fF
C3061 XA6/XA1/XA4/MN1/S AVDD 0.02fF
C3062 XA2/EN EN 1.01fF
C3063 XA3/XA1/XA5/MP2/S AVDD 0.08fF
C3064 XA7/XA1/XA4/MP1/S EN 0.02fF
C3065 XA5/XA2/MP1/a_216_n18# AVDD 0.08fF
C3066 XA8/XA1/XA4/MN2/a_324_n18# XA8/XA1/XA5/MN0/a_324_n18# 0.01fF
C3067 XA0/XA1/XA5/MN2/a_324_n18# XA0/XA1/XA2/Y 0.07fF
C3068 XA2/CN0 SARP 0.02fF
C3069 XA2/XA3/MN2/a_324_n18# AVSS 0.01fF
C3070 XA4/XA2/MP2/a_216_n18# XA4/XA2/MP1/a_216_n18# 0.01fF
C3071 XDAC2/XC1/XRES4/B XDAC2/XC64a<0>/XRES16/B 0.03fF
C3072 XA0/XA9/Y XA0/XA9/MN1/a_324_334# 0.09fF
C3073 XA0/CP0 XA0/XA4/MP1/a_216_n18# 0.02fF
C3074 XA20/XA2/MN6/a_324_n18# XA20/XA3/N1 0.01fF
C3075 XA6/XA7/MN0/a_324_n18# XA6/XA9/B 0.01fF
C3076 XA3/XA7/MP0/a_216_n18# AVDD 0.09fF
C3077 XA6/XA4/A XA5/CN1 0.04fF
C3078 XA3/CN0 D<8> 0.10fF
C3079 XA3/EN XA2/XA1/XA4/MP2/S 0.02fF
C3080 XA4/XA4/A XA4/XA4/MN1/a_324_n18# 0.15fF
C3081 XA2/XA2/A AVDD 1.07fF
C3082 XDAC2/XC64a<0>/XRES4/B XDAC2/XC32a<0>/XRES8/B 0.01fF
C3083 XA7/XA1/XA4/MN2/S XA20/CNO 0.01fF
C3084 XA3/XA1/XA5/MN1/S AVDD 0.02fF
C3085 XA7/XA2/MN3/a_324_n18# XA7/XA2/A 0.15fF
C3086 XA20/XA11/Y DONE 0.06fF
C3087 XB1/XCAPB1/XCAPB0/m3_252_308# XB1/XA4/GNG 0.13fF
C3088 XA3/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C3089 XA0/XA8/MN0/a_324_n18# XA1/EN 0.06fF
C3090 XA0/XA6/MP1/a_216_n18# XA0/CN0 0.15fF
C3091 XA1/XA4/MP2/a_216_n18# AVDD 0.07fF
C3092 XA6/XA11/MP0/a_216_n18# XA6/XA11/MP1/a_216_n18# 0.01fF
C3093 XA3/XA1/XA5/MP1/S AVDD 0.13fF
C3094 XB2/XA3/MP0/S SARN 0.01fF
C3095 XA4/XA9/MN1/a_324_n18# XA4/XA9/A 0.07fF
C3096 XA6/CN1 D<2> 0.42fF
C3097 XA6/XA2/A XA6/XA2/MP1/a_216_n18# 0.15fF
C3098 SARN SARP 6.41fF
C3099 XA20/CNO XA0/XA1/XA1/MN2/S 0.03fF
C3100 XA1/CP0 VREF 0.83fF
C3101 XA4/XA9/A XA3/XA9/A 0.02fF
C3102 XA20/XA3/N2 XA20/XA3/N1 0.51fF
C3103 XA1/XA1/XA4/MP2/S AVDD 0.11fF
C3104 XA2/CN0 XA2/XA6/MP1/S 0.02fF
C3105 XDAC2/XC1/XRES16/B AVDD 0.01fF
C3106 XA8/XA4/MN3/a_324_n18# XA8/CP0 0.02fF
C3107 XA4/XA6/MP1/S CK_SAMPLE 0.03fF
C3108 XA0/XA2/MP2/a_216_n18# AVDD 0.07fF
C3109 XA1/XA1/XA1/MP3/a_216_n18# XA20/CPO 0.08fF
C3110 XA2/XA1/XA5/MP0/a_216_n18# XA2/XA1/XA5/MP1/a_216_n18# 0.01fF
C3111 XA20/XA2a/MN3/a_324_n18# XA20/XA2a/MN2/a_324_n18# 0.01fF
C3112 XDAC2/XC128a<1>/XRES1A/B AVSS 2.97fF
C3113 XA1/XA1/XA1/MP1/a_216_n18# XA1/XA1/XA1/MP3/G 0.01fF
C3114 XA3/EN XA2/XA1/XA1/MP2/a_216_n18# 0.02fF
C3115 AVDD XB1/XA3/MP2/a_216_n18# 0.16fF
C3116 XB2/XA4/MN1/a_324_334# XB2/XA7/MN1/a_324_n18# 0.01fF
C3117 D<0> XA8/XA6/MP2/a_216_n18# 0.07fF
C3118 XA8/XA1/XA1/MP3/a_216_n18# XA8/XA1/XA2/MP0/a_216_n18# 0.01fF
C3119 XA0/XA3/MN2/a_324_n18# D<8> 0.16fF
C3120 XA2/XA1/XA2/MN0/a_324_n18# XA2/XA1/XA4/MN0/a_324_n18# 0.01fF
C3121 XA8/XA1/XA5/MP1/S XA20/CNO 0.03fF
C3122 XA8/EN XA8/XA2/A 0.06fF
C3123 XA0/XA2/MP2/a_216_n18# XA0/XA2/MP1/a_216_n18# 0.01fF
C3124 VREF XA2/CEO 0.32fF
C3125 XA5/XA1/XA1/MN2/S AVSS 0.27fF
C3126 D<5> XA0/CN0 0.05fF
C3127 XA8/XA9/MN0/a_324_n18# XA8/XA9/A 0.15fF
C3128 XDAC2/XC128a<1>/XRES1B/B XDAC2/XC128a<1>/XRES1A/B 0.01fF
C3129 XA2/XA6/MN1/a_324_n18# XA2/XA6/MN2/a_324_n18# 0.01fF
C3130 D<2> XA6/XA3/MP1/a_216_n18# 0.03fF
C3131 XA4/XA3/MP1/a_216_n18# XA4/XA3/MP2/a_216_n18# 0.01fF
C3132 XA5/CP0 XA5/XA5/MP1/a_216_n18# 0.15fF
C3133 XA0/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C3134 XDAC1/XC64a<0>/XRES1B/B AVSS 3.58fF
C3135 XA8/XA3/MP1/a_216_n18# AVDD 0.07fF
C3136 XA20/CPO XA3/XA1/XA2/MN0/a_324_n18# 0.02fF
C3137 XA4/XA2/MN2/a_324_n18# AVSS 0.01fF
C3138 D<1> XA1/CN0 0.04fF
C3139 XA4/XA5/MP3/a_216_n18# XA4/XA5/MP2/a_216_n18# 0.01fF
C3140 XA3/CP0 XA1/CN1 0.04fF
C3141 XA3/XA9/MN1/a_324_334# XA3/XA9/Y 0.09fF
C3142 XA4/XA9/Y AVSS 0.22fF
C3143 XA6/XA4/MP3/a_216_n18# XA6/XA4/MP2/a_216_n18# 0.01fF
C3144 XB2/XA4/MN1/S XB2/XA4/GNG 0.01fF
C3145 XDAC2/XC64b<1>/XRES16/B XDAC2/X16ab/XRES16/B 0.41fF
C3146 XA0/XA5/MP1/a_216_n18# XA0/XA5/MP2/a_216_n18# 0.01fF
C3147 XDAC1/XC1/XRES8/B SARP 11.94fF
C3148 XA4/XA1/XA1/MP3/S AVSS 0.02fF
C3149 XA1/XA1/XA5/MN2/a_324_n18# XA1/XA1/XA5/MN1/a_324_n18# 0.01fF
C3150 XA20/XA3/MN4/a_324_n18# SARN 0.15fF
C3151 XA6/XA2/MN0/a_324_n18# AVSS 0.01fF
C3152 XA5/XA5/MN3/a_324_n18# XA5/XA5/MN2/a_324_n18# 0.01fF
C3153 XA7/XA2/MP1/a_216_n18# XA7/XA2/MP2/a_216_n18# 0.01fF
C3154 XA6/XA1/XA5/MP2/S VREF 0.03fF
C3155 XDAC1/X16ab/XRES16/B AVSS 16.03fF
C3156 XA4/XA1/XA4/MN2/S XA20/CNO 0.01fF
C3157 XA8/XA4/MP0/a_216_n18# AVDD 0.08fF
C3158 XDAC2/XC64b<1>/XRES1A/B XDAC2/XC0/XRES1A/B 0.03fF
C3159 XA6/XA1/XA2/Y XA6/XA1/XA5/MN0/a_324_n18# 0.02fF
C3160 XDAC2/XC64b<1>/XRES1A/B XDAC2/XC64b<1>/XRES8/B 0.12fF
C3161 XDAC2/XC64b<1>/XRES2/B XDAC2/XC64b<1>/XRES4/B 0.55fF
C3162 XA1/XA1/XA2/Y XA20/CNO 0.22fF
C3163 XA1/XA1/XA5/MP1/S XA20/CNO 0.01fF
C3164 XA8/XA5/MN2/a_324_n18# XA8/XA5/MN1/a_324_n18# 0.01fF
C3165 XA20/XA10/MN1/a_324_n18# XA20/XA11/Y 0.08fF
C3166 XA6/XA12/MN0/a_324_n18# XA6/XA12/A 0.09fF
C3167 XDAC2/XC128b<2>/XRES4/B XDAC2/X16ab/XRES1A/B 0.01fF
C3168 XDAC1/X16ab/XRES1B/B XDAC1/X16ab/XRES16/B 0.12fF
C3169 XA3/XA1/XA1/MN0/a_324_n18# XA3/XA1/XA1/MN1/a_324_n18# 0.01fF
C3170 D<0> XA8/XA2/A 0.02fF
C3171 XA4/XA11/MN1/a_324_n18# AVSS 0.01fF
C3172 XA3/XA1/XA0/MN1/a_324_n18# XA3/XA1/XA1/MN0/a_324_n18# 0.01fF
C3173 XDAC2/XC128a<1>/XRES16/B XDAC2/XC32a<0>/XRES2/B 0.01fF
C3174 XA3/XA4/MP3/a_216_n18# XA3/XA5/MP0/a_216_n18# 0.01fF
C3175 XA3/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C3176 XDAC1/XC1/XRES4/B AVSS 5.45fF
C3177 XA8/ENO XA8/XA1/XA4/MP0/a_216_n18# 0.08fF
C3178 AVDD XA2/XA1/XA1/MP1/a_216_n18# 0.08fF
C3179 XA3/XA11/A XA3/XA12/A 0.07fF
C3180 XA8/XA9/B XA8/XA9/Y 0.15fF
C3181 XA7/XA1/XA4/MN1/S XA20/CPO 0.04fF
C3182 SARN XA20/XA4/MN4/a_324_n18# 0.15fF
C3183 XA2/XA9/B XA2/XA6/MP3/S 0.07fF
C3184 XA5/EN XA5/XA1/XA2/Y 0.14fF
C3185 XA7/XA12/A XA7/XA13/MP1/a_216_n18# 0.08fF
C3186 XB2/XA3/MN2/a_324_n18# XB2/XA4/MN0/a_324_n18# 0.01fF
C3187 XA3/XA9/MP1/a_216_n18# XA3/XA9/MP0/a_216_n18# 0.01fF
C3188 XA0/XA5/MP2/a_216_n18# AVDD 0.07fF
C3189 XA6/CN0 XA6/XA6/MP2/a_216_n18# 0.08fF
C3190 XA5/XA1/XA4/MN1/S AVDD 0.02fF
C3191 XA8/XA13/MN1/a_324_334# XA8/XA13/MN1/a_324_n18# 0.01fF
C3192 XA2/XA1/XA1/MP2/S XA3/EN 0.14fF
C3193 XA7/XA9/A XA8/XA9/B 0.02fF
C3194 XA1/XA1/XA1/MP3/S XA20/CPO 0.01fF
C3195 XA2/XA1/XA1/MP3/G AVSS 0.12fF
C3196 XA8/ENO XA8/XA1/XA1/MP3/G 0.24fF
C3197 XA8/XA9/MP0/a_216_n18# AVDD 0.09fF
C3198 XA6/XA5/MN2/a_324_n18# AVSS 0.01fF
C3199 XA7/XA2/MN1/a_324_n18# XA7/XA2/MN0/a_324_n18# 0.01fF
C3200 XA1/XA3/MP1/a_216_n18# XA1/XA3/MP2/a_216_n18# 0.01fF
C3201 AVDD XA0/XA1/XA1/MP1/a_216_n18# 0.08fF
C3202 XA8/EN XA7/XA1/XA1/MP3/a_216_n18# 0.01fF
C3203 XA3/CN1 XA1/CN0 0.20fF
C3204 XA3/XA11/MN0/a_324_n18# XA3/XA9/Y 0.07fF
C3205 XA0/XA11/MN1/a_324_n18# XA0/XA11/MN0/a_324_n18# 0.01fF
C3206 XA7/XA9/MP1/a_216_n18# XA7/XA9/A 0.08fF
C3207 XA4/CN0 XA4/EN 0.03fF
C3208 XA1/CN0 XA1/XA5/MP2/a_216_n18# 0.01fF
C3209 XA6/CN1 XA8/EN 0.03fF
C3210 XA5/CP0 XA5/XA5/MN0/a_324_n18# 0.09fF
C3211 XA0/XA12/A XA0/XA13/MP1/a_216_n18# 0.08fF
C3212 XA8/XA1/XA5/MN1/S XA20/CNO 0.03fF
C3213 XA6/XA9/MP0/a_216_n18# XA6/XA8/MP0/a_216_n18# 0.01fF
C3214 XA6/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C3215 XA20/XA2/MP5/a_216_n18# XA20/XA2/MP6/a_216_n18# 0.01fF
C3216 XA3/XA1/XA5/MN2/a_324_n18# XA3/XA1/XA2/Y 0.07fF
C3217 XA3/CP0 XA3/XA1/XA1/MP3/G 0.02fF
C3218 XA6/XA4/MP3/a_216_n18# XA6/CP0 0.02fF
C3219 XA20/CNO XA0/XA1/XA1/MP3/G 0.06fF
C3220 XA7/XA6/MP1/S AVDD 0.12fF
C3221 XA6/XA1/XA4/MP2/S XA7/EN 0.02fF
C3222 AVDD XB1/XA3/MP0/a_216_n18# 0.08fF
C3223 XA4/XA5/MP2/a_216_n18# XA4/CN0 0.01fF
C3224 XA7/XA1/XA1/MN1/a_324_n18# AVSS 0.01fF
C3225 XA20/XA9/Y XA20/XA3/MP4/a_216_n18# 0.08fF
C3226 XA0/XA9/Y XA0/XA11/MN0/a_324_n18# 0.07fF
C3227 SAR_IN XB2/M3/a_324_n18# 0.02fF
C3228 XA20/XA4/MN3/a_324_n18# XA20/XA4/MN4/a_324_n18# 0.01fF
C3229 XA3/XA1/XA2/Y AVDD 0.33fF
C3230 XA2/CN0 XDAC2/X16ab/XRES16/B 0.03fF
C3231 XA7/XA9/B XA7/XA8/MN0/a_324_n18# 0.01fF
C3232 XA5/XA4/MP1/a_216_n18# AVDD 0.07fF
C3233 D<2> XA1/CN0 0.07fF
C3234 XA6/XA5/MP1/a_216_n18# AVDD 0.07fF
C3235 SARN XB1/M7/a_324_n18# 0.02fF
C3236 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC0/XRES16/B 0.05fF
C3237 XB1/XA3/B XB1/XA5b/MP1/a_216_n18# 0.02fF
C3238 AVDD XA2/XA1/XA4/MP2/a_216_n18# 0.08fF
C3239 XA2/XA1/XA5/MP2/a_216_n18# XA2/XA1/XA5/MP1/a_216_n18# 0.01fF
C3240 XA20/XA9/Y SARP 0.43fF
C3241 XA4/XA6/MN0/a_324_n18# XA4/CP0 0.07fF
C3242 XB2/XA1/Y XB2/M4/G 0.12fF
C3243 XA2/XA6/MP3/a_216_n18# D<6> 0.15fF
C3244 XA8/XA1/XA4/MP2/S XA20/CNO 0.01fF
C3245 XA5/CP0 XA6/EN 0.06fF
C3246 XA2/XA1/XA5/MN1/a_324_n18# XA2/XA1/XA5/MN2/a_324_n18# 0.01fF
C3247 XA6/XA4/A XA7/EN 0.11fF
C3248 XA0/XA1/XA4/MN2/S AVDD 0.02fF
C3249 XA7/CN0 XA1/CN0 0.12fF
C3250 XA2/CN0 XA4/CN0 0.08fF
C3251 XA7/XA5/MN3/a_324_n18# XA7/CP0 0.15fF
C3252 XA1/XA2/A XA1/EN 0.09fF
C3253 XA20/CPO XA3/XA1/XA1/MP3/a_216_n18# 0.08fF
C3254 XA3/XA4/MN0/a_324_n18# AVSS 0.01fF
C3255 XA6/XA11/MP1/S AVDD 0.19fF
C3256 D<5> D<6> 0.24fF
C3257 XA1/XA4/A XA1/XA4/MN0/a_324_n18# 0.09fF
C3258 XA20/CNO D<8> 0.15fF
C3259 XA0/CP1 XA0/XA9/B 0.05fF
C3260 CK_SAMPLE_BSSW XB1/XA0/MP0/a_216_n18# 0.07fF
C3261 XA4/XA1/XA2/Y XA3/XA1/XA2/Y 0.02fF
C3262 XA2/CN0 XA5/CN0 0.09fF
C3263 XDAC2/X16ab/XRES16/B SARN 21.64fF
C3264 VREF XA2/XA1/XA5/MP1/S 0.02fF
C3265 XA1/XA2/MN3/a_324_n18# XA1/XA2/MN2/a_324_n18# 0.01fF
C3266 D<3> XA1/CN0 0.12fF
C3267 XA4/XA1/XA5/MP0/a_216_n18# XA4/XA1/XA5/MP1/a_216_n18# 0.01fF
C3268 XA2/XA4/A XA20/CNO 0.18fF
C3269 XA3/CN1 XA3/EN 0.22fF
C3270 XA0/XA3/MP3/a_216_n18# AVDD 0.07fF
C3271 VREF XA8/XA9/Y 0.02fF
C3272 XA0/XA3/MP2/a_216_n18# AVDD 0.07fF
C3273 XA20/XA3/MP3/a_216_n18# AVDD 0.17fF
C3274 XA8/XA9/MN1/a_324_334# XA8/XA9/MN1/a_324_n18# 0.01fF
C3275 XDAC1/XC64b<1>/XRES8/B XDAC1/XC0/XRES16/B 0.03fF
C3276 AVSS XA3/XA4/A 1.07fF
C3277 XB1/XCAPB1/XCAPB2/m3_9756_132# XB1/XA4/GNG 0.02fF
C3278 XA3/CEO XA4/XA12/A 0.14fF
C3279 XDAC1/XC32a<0>/XRES16/B XDAC1/XC32a<0>/XRES2/B 1.61fF
C3280 XA4/XA1/XA2/MN0/a_324_n18# XA20/CPO 0.01fF
C3281 XA4/CN0 SARN 0.07fF
C3282 XA1/XA1/XA4/MN1/S XA20/CPO 0.04fF
C3283 XA0/CEO AVSS 0.49fF
C3284 XA20/XA9/A SARP 0.40fF
C3285 XA7/XA9/A VREF 0.04fF
C3286 XB2/XA5/MP1/a_216_334# AVDD 0.17fF
C3287 XA2/XA7/MN0/a_324_n18# XA2/XA6/MN3/a_324_n18# 0.01fF
C3288 XA0/XA1/XA4/MP1/a_216_n18# XA0/XA1/XA4/MP2/a_216_n18# 0.01fF
C3289 XA7/XA3/MN2/a_324_n18# XA7/XA3/MN1/a_324_n18# 0.01fF
C3290 XA6/CN0 AVSS 1.00fF
C3291 XA2/XA9/MN0/a_324_n18# XA2/XA8/MN0/a_324_n18# 0.01fF
C3292 D<0> XA8/XA6/MP1/S 0.02fF
C3293 XA20/XA2/MN4/a_324_n18# SARP 0.15fF
C3294 XA5/XA1/XA1/MP2/a_216_n18# XA20/CPO 0.06fF
C3295 XA5/CN0 SARN 0.07fF
C3296 XA20/CPO XA0/XA1/XA4/MN1/a_324_n18# 0.07fF
C3297 XA0/XA1/XA5/MP1/a_216_n18# XA0/XA1/XA5/MP2/a_216_n18# 0.01fF
C3298 XA5/XA1/XA4/MP1/S AVDD 0.14fF
C3299 XA7/XA4/A AVDD 1.42fF
C3300 XA7/XA13/MP1/a_216_334# AVDD 0.17fF
C3301 XA3/XA1/XA4/MP1/S XA3/XA1/XA4/MP2/S 0.04fF
C3302 AVDD XA2/XA11/MP1/a_216_n18# 0.08fF
C3303 EN XA2/XA1/XA1/MP3/G 0.10fF
C3304 XA3/XA5/MN0/a_324_n18# XA3/XA4/A 0.07fF
C3305 XB2/XA2/MP0/G XA0/CEIN 0.04fF
C3306 AVDD XA2/XA1/XA5/MP1/a_216_n18# 0.08fF
C3307 XA3/XA5/MP1/a_216_n18# VREF 0.02fF
C3308 D<5> SARP 0.16fF
C3309 XA6/XA1/XA2/Y AVSS 0.31fF
C3310 XA1/XA12/A AVDD 0.44fF
C3311 XB1/XA2/MP0/G XB1/XA1/Y 0.01fF
C3312 XDAC1/XC1/XRES2/B XDAC1/XC64a<0>/XRES2/B 0.05fF
C3313 XA8/XA6/MP2/a_216_n18# XA8/CN0 0.08fF
C3314 XA3/XA1/XA4/MN2/S AVDD 0.02fF
C3315 XA3/XA6/MN3/a_324_n18# XA3/XA6/MN2/a_324_n18# 0.01fF
C3316 XA0/XA5/MP1/a_216_n18# XA0/CN0 0.02fF
C3317 XA3/CEO XA4/XA12/MN0/a_324_n18# 0.07fF
C3318 XA4/XA9/Y XA4/XA9/A 0.04fF
C3319 XA6/XA1/XA5/MP2/a_216_n18# EN 0.16fF
C3320 XA5/XA2/A AVDD 1.07fF
C3321 XA2/EN XA2/CN1 0.22fF
C3322 XA6/XA3/MP0/a_216_n18# XA6/CN1 0.07fF
C3323 XA4/XA2/MP1/a_216_n18# VREF 0.02fF
C3324 XA3/XA11/MP1/S AVDD 0.18fF
C3325 XA20/XA2/MN1/a_324_n18# XA20/XA9/Y 0.07fF
C3326 XA8/ENO XA8/XA2/A 0.10fF
C3327 XA2/XA3/MP0/a_216_n18# XA2/XA2/A 0.08fF
C3328 XA5/EN XA5/XA1/XA4/MN1/S 0.02fF
C3329 XA1/XA1/XA2/Y XA2/XA1/XA2/Y 0.02fF
C3330 XA3/XA1/XA5/MP2/a_216_n18# XA3/XA1/XA5/MP1/a_216_n18# 0.01fF
C3331 XDAC1/XC1/XRES16/B XDAC1/XC64a<0>/XRES1A/B 0.04fF
C3332 XA2/CP0 XA2/XA4/MP1/a_216_n18# 0.02fF
C3333 XA8/XA1/XA5/MN1/S XA8/XA1/XA5/MN2/S 0.04fF
C3334 XA2/CN0 XA2/XA5/MP2/a_216_n18# 0.01fF
C3335 XA0/XA5/MN3/a_324_n18# XA0/CN0 0.01fF
C3336 XB2/XCAPB1/XCAPB2/m3_324_308# XB2/XA4/GNG 0.07fF
C3337 XA3/CEO XA4/XA11/A 0.08fF
C3338 XA6/EN XA20/CNO 1.02fF
C3339 XA1/XA2/A XA2/XA2/A 0.03fF
C3340 XA1/XA13/MP1/a_216_334# AVDD 0.17fF
C3341 XA6/XA3/MP0/a_216_n18# XA6/XA3/MP1/a_216_n18# 0.01fF
C3342 XA8/ENO XA8/XA1/XA4/MP1/S 0.02fF
C3343 XB1/XA7/MN1/a_324_334# XB1/XA7/MN1/a_324_n18# 0.01fF
C3344 XA6/XA6/MP3/S AVDD 0.16fF
C3345 XA20/XA1/MN0/a_324_n18# XA20/XA0/MN1/a_324_n18# 0.01fF
C3346 XA3/XA4/MN0/a_324_n18# XA3/XA3/MN3/a_324_n18# 0.01fF
C3347 XDAC1/XC0/XRES1A/B XDAC1/XC0/XRES16/B 1.60fF
C3348 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC0/XRES1B/B 0.03fF
C3349 XA8/XA2/MP2/a_216_n18# VREF 0.03fF
C3350 XA6/XA1/XA1/MP2/a_216_n18# XA20/CPO 0.06fF
C3351 XA5/CEO XA6/XA12/A 0.14fF
C3352 XA2/XA12/A XA2/XA13/MP1/a_216_n18# 0.08fF
C3353 AVDD XA0/CN0 5.57fF
C3354 XA7/XA6/MP2/a_216_n18# AVDD 0.09fF
C3355 XA6/XA9/B XA6/XA8/MN0/a_324_n18# 0.01fF
C3356 D<1> XA7/XA3/MP3/a_216_n18# 0.02fF
C3357 XA6/CN0 CK_SAMPLE 0.07fF
C3358 XA7/XA1/XA1/MP2/S XA7/XA1/XA1/MP3/G 0.04fF
C3359 XA4/XA1/XA5/MP1/S EN 0.03fF
C3360 XA20/XA11/MP1/S AVDD 0.17fF
C3361 XB2/XA3/B XB2/XCAPB1/XCAPB1/m3_9828_132# 0.21fF
C3362 XA5/XA9/B XA5/XA8/MN0/a_324_n18# 0.01fF
C3363 XA1/XA9/MN1/a_324_n18# XA1/XA9/A 0.07fF
C3364 VREF XA0/XA12/A 0.03fF
C3365 XDAC1/XC32a<0>/XRES8/B XDAC1/XC128a<1>/XRES8/B 0.21fF
C3366 EN XA3/XA4/A 0.09fF
C3367 XDAC2/XC1/XRES8/B SARN 11.94fF
C3368 XA6/XA5/MP0/a_216_n18# XA6/XA5/MP1/a_216_n18# 0.01fF
C3369 XDAC1/XC64b<1>/XRES4/B XDAC1/XC64b<1>/XRES1A/B 0.29fF
C3370 XA3/XA3/MN3/a_324_n18# XA3/XA4/A 0.01fF
C3371 XA20/XA3/N1 XA20/CPO 0.25fF
C3372 XA1/XA9/MP0/a_216_n18# AVDD 0.09fF
C3373 XA1/XA13/MP1/a_216_n18# AVDD 0.13fF
C3374 XA3/CP0 AVSS 1.32fF
C3375 XA3/CEO XA3/XA12/A 0.20fF
C3376 XB1/XA3/MP0/a_216_334# XB1/XA3/MP2/a_216_n18# 0.01fF
C3377 XA6/CN0 EN 0.07fF
C3378 XA20/XA12/MN0/a_324_n18# AVSS 0.01fF
C3379 XA0/XA11/MN1/a_324_n18# XA0/CEIN 0.08fF
C3380 XA3/XA13/MN1/a_324_n18# AVSS 0.09fF
C3381 XDAC1/XC64b<1>/XRES1B/B SARP 1.79fF
C3382 XA8/XA1/XA4/MN2/S XA20/CPO 0.01fF
C3383 XA6/XA4/A XA6/XA4/MP2/a_216_n18# 0.15fF
C3384 XA6/XA9/MN1/a_324_n18# XA6/XA9/MN0/a_324_n18# 0.01fF
C3385 XB2/XA1/Y XB2/XA1/MP0/G 0.13fF
C3386 XA8/XA6/MN0/a_324_n18# XA8/CP0 0.07fF
C3387 XDAC1/X16ab/XRES1A/B XDAC1/X16ab/XRES16/B 1.60fF
C3388 XA0/XA1/XA5/MN2/S XA20/CNO 0.01fF
C3389 XA1/EN XA1/CN1 0.21fF
C3390 XDAC1/XC128a<1>/XRES16/B XDAC1/XC128a<1>/XRES1A/B 1.60fF
C3391 XA2/XA5/MP3/a_216_n18# XA2/XA5/MP2/a_216_n18# 0.01fF
C3392 XA0/XA5/MN1/a_324_n18# XA0/XA5/MN2/a_324_n18# 0.01fF
C3393 XA2/EN D<7> 0.46fF
C3394 XA0/XA9/Y XA0/CEIN 0.01fF
C3395 XA2/XA5/MP1/a_216_n18# XA2/XA5/MP0/a_216_n18# 0.01fF
C3396 XA0/XA3/MN3/a_324_n18# XA0/XA3/MN2/a_324_n18# 0.01fF
C3397 XA4/XA9/MP1/a_216_n18# XA4/XA9/A 0.08fF
C3398 XA1/XA9/MP1/a_216_334# AVDD 0.09fF
C3399 XDAC2/XC1/XRES1B/B XDAC2/XC1/XRES8/B 0.12fF
C3400 XA8/EN XA8/XA1/XA1/MN1/a_324_n18# 0.08fF
C3401 XDAC1/XC32a<0>/XRES1B/B SARP 1.79fF
C3402 XA2/XA1/XA1/MN0/a_324_n18# XA2/XA1/XA1/MN1/a_324_n18# 0.01fF
C3403 XA0/XA1/XA4/MN2/a_324_n18# XA0/XA1/XA4/MN1/a_324_n18# 0.01fF
C3404 XA7/XA2/MN2/a_324_n18# XA7/XA2/MN3/a_324_n18# 0.01fF
C3405 D<7> XA1/XA6/MP3/a_216_n18# 0.15fF
C3406 XA20/XA3/MP3/a_216_n18# XA20/XA3/MP2/a_216_n18# 0.01fF
C3407 XA4/XA1/XA4/MN2/S XA4/XA1/XA4/MP2/S 0.01fF
C3408 XA6/XA1/XA2/Y EN 0.07fF
C3409 XA2/XA3/MP3/a_216_n18# AVDD 0.07fF
C3410 XA8/XA1/XA1/MP3/S AVDD 0.14fF
C3411 XA6/XA1/XA4/MN2/a_324_n18# XA6/XA1/XA5/MN0/a_324_n18# 0.01fF
C3412 XA3/CP0 XA3/XA5/MN0/a_324_n18# 0.09fF
C3413 XA2/XA4/A XA2/XA5/MP0/a_216_n18# 0.08fF
C3414 XA4/XA8/MP0/a_216_n18# XA4/XA7/MP0/a_216_n18# 0.01fF
C3415 XA1/XA1/XA1/MN0/a_324_n18# XA1/EN 0.09fF
C3416 XA6/XA2/MN0/a_324_n18# XA6/XA2/MN1/a_324_n18# 0.01fF
C3417 XDAC2/XC0/XRES1B/B XDAC2/XC0/XRES16/B 0.13fF
C3418 XB2/CKN XA0/CEIN 0.08fF
C3419 XA6/CN1 XA7/CN1 0.03fF
C3420 XDAC1/XC128b<2>/XRES8/B XDAC1/X16ab/XRES16/B 0.03fF
C3421 XA7/CEO XA8/XA12/A 0.14fF
C3422 XA6/XA1/XA5/MP1/S XA6/XA1/XA5/MN1/S 0.01fF
C3423 XA5/XA1/XA5/MP1/S AVDD 0.13fF
C3424 XA3/XA5/MN3/a_324_n18# XA3/XA6/MN0/a_324_n18# 0.01fF
C3425 XA8/XA3/MN1/a_324_n18# XA8/CN1 0.16fF
C3426 XDAC2/XC128b<2>/XRES1B/B XDAC2/X16ab/XRES16/B 0.05fF
C3427 XDAC1/XC128a<1>/XRES1B/B SARP 1.79fF
C3428 XA0/XA5/MP3/a_216_n18# AVDD 0.07fF
C3429 XA2/CN1 XA2/XA3/MN2/a_324_n18# 0.16fF
C3430 XA3/XA5/MP3/a_216_n18# AVDD 0.07fF
C3431 XA2/XA4/A XA2/XA1/XA2/Y 0.19fF
C3432 XDAC2/XC1/XRES16/B XDAC2/XC1/XRES1A/B 1.61fF
C3433 XA0/CP0 D<4> 0.10fF
C3434 XA0/CP1 XA20/CNO 0.05fF
C3435 XA6/XA9/B VREF 0.12fF
C3436 XDAC2/XC128a<1>/XRES8/B SARN 11.94fF
C3437 XA5/CN1 AVDD 1.31fF
C3438 XDAC2/XC128a<1>/XRES16/B XDAC2/XC32a<0>/XRES16/B 0.41fF
C3439 XDAC2/XC64b<1>/XRES2/B XDAC2/X16ab/XRES2/B 0.05fF
C3440 XA0/XA8/MN0/a_324_n18# XA0/XA7/MN0/a_324_n18# 0.01fF
C3441 XA3/XA1/XA4/MP0/a_216_n18# XA4/EN 0.08fF
C3442 XA1/CP0 XDAC1/XC64b<1>/XRES16/B 0.01fF
C3443 XA3/CN0 XA4/EN 0.15fF
C3444 XA3/XA2/MN0/a_324_n18# XA3/EN 0.07fF
C3445 XA0/XA9/Y XA0/XA9/MP1/a_216_334# 0.07fF
C3446 XA4/XA5/MP3/a_216_n18# XA4/CP0 0.15fF
C3447 XA2/DONE AVDD 0.21fF
C3448 AVDD XA1/XA5/MP1/a_216_n18# 0.07fF
C3449 XA6/XA1/XA2/MN0/a_324_n18# XA20/CPO 0.01fF
C3450 XB2/XCAPB1/XCAPB3/m3_9756_132# XB2/XA4/GNG 0.02fF
C3451 XA0/XA1/XA2/MP0/a_216_n18# XA1/EN 0.08fF
C3452 XA5/XA2/A XA5/EN 0.09fF
C3453 XA1/EN XA0/XA1/XA1/MP0/a_216_n18# 0.01fF
C3454 XA3/XA9/A VREF 0.04fF
C3455 XA8/XA9/A XA8/XA9/Y 0.04fF
C3456 XDAC1/XC32a<0>/XRES16/B XA1/CP0 0.02fF
C3457 EN XA0/XA1/XA5/MP2/S 0.04fF
C3458 XA0/CP1 XA0/XA6/MP3/a_216_n18# 0.15fF
C3459 XA4/DONE AVDD 0.21fF
C3460 XA1/XA4/MN0/a_324_n18# XA1/XA3/MN3/a_324_n18# 0.01fF
C3461 XA6/EN XA5/XA9/A 0.09fF
C3462 XA20/XA1/MP3_DMY/a_216_n18# XA20/XA1/MP2_DMY/a_216_n18# 0.01fF
C3463 XA0/XA13/MP1/a_216_n18# XA0/XA13/MP1/a_216_334# 0.01fF
C3464 XA4/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C3465 XA6/XA4/A XA6/CP0 0.52fF
C3466 XA20/XA9/Y DONE 0.02fF
C3467 XA7/XA12/A XA7/XA12/MN0/a_324_n18# 0.09fF
C3468 XA0/XA1/XA4/MP1/S AVDD 0.14fF
C3469 XA3/CP0 CK_SAMPLE 0.09fF
C3470 XA7/XA9/A XA8/XA9/A 0.02fF
C3471 XA3/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C3472 XA0/XA2/A VREF 0.36fF
C3473 XA3/CN0 XA2/CN0 0.55fF
C3474 AVDD XA3/XA4/MP3/a_216_n18# 0.07fF
C3475 XA8/CN0 XA8/XA5/MN1/a_324_n18# 0.02fF
C3476 XA2/CP0 XA0/CP0 0.42fF
C3477 XA1/XA4/A XA1/XA4/MP1/a_216_n18# 0.15fF
C3478 XA20/CPO XA0/XA1/XA1/MP2/a_216_n18# 0.06fF
C3479 XB2/XA3/MP0/S XB2/XA4/MN0/a_324_n18# 0.07fF
C3480 XA20/XA2/N2 XA20/XA3a/A 0.14fF
C3481 XA1/XA1/XA1/MN2/S D<7> 0.01fF
C3482 XA6/XA7/MP0/a_216_n18# XA6/XA8/MP0/a_216_n18# 0.01fF
C3483 XA7/XA1/XA2/MN0/a_324_n18# XA20/CPO 0.02fF
C3484 XA2/EN VREF 1.22fF
C3485 XA6/XA1/XA5/MP2/a_216_n18# XA6/XA1/XA5/MP1/a_216_n18# 0.01fF
C3486 XA2/XA9/MP1/a_216_n18# XA2/XA9/B 0.07fF
C3487 XA8/XA1/XA5/MP1/S XA8/XA4/A 0.02fF
C3488 XA8/XA1/XA1/MP2/a_216_n18# XA20/CNO 0.08fF
C3489 XA1/XA1/XA1/MP3/G XA1/CN0 0.02fF
C3490 XA5/XA9/Y AVDD 0.58fF
C3491 XA8/CEO XA8/XA13/MP1/a_216_n18# 0.01fF
C3492 XA3/CP0 EN 0.05fF
C3493 XA8/CN0 XA8/XA6/MP1/S 0.02fF
C3494 XA20/XA2/MN2/a_324_n18# XA20/XA2/N2 0.01fF
C3495 XA3/XA9/MN1/a_324_334# XA3/XA9/B 0.07fF
C3496 D<6> AVDD 1.85fF
C3497 XA5/XA1/XA1/MP2/S XA5/XA1/XA1/MP3/S 0.04fF
C3498 XA2/XA2/A XA1/CN1 0.03fF
C3499 XA0/XA4/A AVDD 1.42fF
C3500 XA2/XA6/MN0/a_324_n18# AVSS 0.01fF
C3501 XB1/XA3/MP0/a_216_334# XB1/XA3/MP0/a_216_n18# 0.01fF
C3502 XA7/XA5/MP3/a_216_n18# XA7/CP0 0.15fF
C3503 XA3/CN0 SARN 0.07fF
C3504 XA6/XA12/A XA6/XA13/MP1/a_216_n18# 0.08fF
C3505 XA1/XA1/XA1/MN1/a_324_n18# XA20/CNO 0.07fF
C3506 XA7/XA4/A XA7/XA2/A 0.14fF
C3507 SARP XB1/M4/G 0.24fF
C3508 XA20/XA11/MN0/a_324_n18# XA20/XA11/Y 0.02fF
C3509 XA20/XA9/A DONE 0.08fF
C3510 XA20/CNO XA2/XA1/XA5/MN2/S 0.01fF
C3511 XA5/XA11/A AVDD 0.45fF
C3512 D<5> XA3/XA3/MP2/a_216_n18# 0.01fF
C3513 XB1/CKN XB1/XA3/MP2/a_216_n18# 0.07fF
C3514 XB2/XCAPB1/XCAPB3/m3_252_308# XB2/XA3/B 0.02fF
C3515 D<4> XA4/XA4/A 0.26fF
C3516 XA6/CN1 XA6/XA4/MN0/a_324_n18# 0.07fF
C3517 XA1/CP0 XA20/CPO 0.06fF
C3518 XA5/EN XA5/XA1/XA5/MN2/a_324_n18# 0.08fF
C3519 XA3/XA1/XA4/MP2/S AVDD 0.11fF
C3520 XB1/XCAPB1/XCAPB1/m3_9828_132# XB1/XA3/B 0.21fF
C3521 AVDD XA20/XA2a/MP3/a_216_n18# 0.09fF
C3522 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MN2/S 0.08fF
C3523 XA7/XA6/MN1/S XA7/XA9/B 0.05fF
C3524 XA6/XA3/MP2/a_216_n18# XA6/CN1 0.15fF
C3525 XA3/XA13/MP1/a_216_n18# XA3/XA12/A 0.08fF
C3526 XDAC1/XC1/XRES1B/B XDAC1/XC1/XRES2/B 0.23fF
C3527 XA4/CN0 XA4/CP0 0.59fF
C3528 XA0/XA9/MN1/S AVSS 0.15fF
C3529 XDAC2/XC64a<0>/XRES1A/B XDAC2/XC64a<0>/XRES4/B 0.29fF
C3530 XA20/CNO XA2/XA1/XA5/MN0/a_324_n18# 0.09fF
C3531 XA2/EN XA2/XA1/XA1/MN0/a_324_n18# 0.08fF
C3532 XA1/XA9/MP0/a_216_n18# XA1/XA9/A 0.14fF
C3533 VREF XA8/XA5/MP2/a_216_n18# 0.03fF
C3534 XA6/XA1/XA4/MP0/a_216_n18# EN 0.07fF
C3535 XA0/XA9/A XA0/XA11/A 0.01fF
C3536 XA20/XA3/MP4/a_216_n18# AVDD 0.09fF
C3537 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC64a<0>/XRES8/B 0.12fF
C3538 XB2/XA3/MP0/S AVDD 0.23fF
C3539 XA20/XA3/CO AVSS 0.31fF
C3540 XA8/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C3541 XA4/XA2/A XA4/XA2/MP1/a_216_n18# 0.15fF
C3542 XA5/XA1/XA5/MN1/S AVSS 0.12fF
C3543 XA4/XA1/XA5/MP2/S EN 0.04fF
C3544 XDAC1/XC64b<1>/XRES4/B XDAC1/XC64b<1>/XRES2/B 0.55fF
C3545 XA2/XA1/XA0/MP1/a_216_n18# XA2/XA1/XA1/MP0/a_216_n18# 0.01fF
C3546 AVDD SARP 0.60fF
C3547 XA4/XA6/MP1/S VREF 0.04fF
C3548 XA0/XA4/MP2/a_216_n18# VREF 0.03fF
C3549 XA6/XA6/MN0/a_324_n18# AVSS 0.01fF
C3550 XA6/XA3/MP2/a_216_n18# XA6/XA3/MP1/a_216_n18# 0.01fF
C3551 XA0/XA1/XA5/MP1/S XA0/XA1/XA5/MN1/S 0.01fF
C3552 XA1/XA1/XA4/MP1/a_216_n18# XA1/XA1/XA4/MP0/a_216_n18# 0.01fF
C3553 XB1/CKN XB1/XA3/MN2/a_324_n18# 0.07fF
C3554 XA0/XA11/MP1/a_216_n18# AVDD 0.08fF
C3555 XB2/XA4/MP1/a_216_334# XB2/XA4/MP1/a_216_n18# 0.01fF
C3556 XA1/XA11/A XA1/CEO 0.05fF
C3557 XA2/CN1 XA2/XA1/XA1/MP3/G 0.02fF
C3558 XDAC1/XC128b<2>/XRES16/B SARP 21.64fF
C3559 XA3/XA11/MN1/a_324_n18# AVSS 0.01fF
C3560 XB1/XA2/MP0/G AVSS 0.09fF
C3561 XDAC1/XC64a<0>/XRES16/B AVSS 16.06fF
C3562 XDAC1/XC1/XRES1A/B XDAC1/XC64a<0>/XRES1A/B 0.03fF
C3563 XDAC2/XC64a<0>/XRES16/B SARN 21.64fF
C3564 XA6/XA4/MN1/a_324_n18# XA6/CP0 0.03fF
C3565 XA2/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C3566 XA3/XA3/MN1/a_324_n18# XA3/CN1 0.16fF
C3567 XA5/CN1 XA5/EN 0.04fF
C3568 XA2/CP0 XA2/XA5/MN0/a_324_n18# 0.09fF
C3569 XA0/XA6/MN3/S AVDD 0.01fF
C3570 AVDD XA2/XA11/MP0/a_216_n18# 0.09fF
C3571 AVDD XA1/XA5/MP3/a_216_n18# 0.07fF
C3572 XA8/XA2/MP3/a_216_n18# AVDD 0.07fF
C3573 XA8/XA1/XA5/MN1/S XA8/XA4/A 0.02fF
C3574 XA2/XA6/MP1/S AVDD 0.12fF
C3575 XA7/XA9/MP1/a_216_n18# XA7/XA9/MP0/a_216_n18# 0.01fF
C3576 XA0/CP0 XA0/XA4/MN3/a_324_n18# 0.02fF
C3577 XA0/XA11/MN1/a_324_n18# XA0/XA12/MN0/a_324_n18# 0.01fF
C3578 XA0/XA3/MP0/a_216_n18# XA0/XA2/A 0.08fF
C3579 XDAC2/XC128b<2>/XRES2/B AVSS 3.71fF
C3580 D<3> XA5/XA4/MP0/a_216_n18# 0.01fF
C3581 XA6/CN0 XA6/XA1/XA1/MP3/G 0.02fF
C3582 XA0/CN0 XDAC2/XC32a<0>/XRES16/B 0.05fF
C3583 XA2/XA9/MN0/a_324_n18# XA2/XA9/B 0.01fF
C3584 XA4/XA1/XA5/MP0/a_216_n18# XA4/XA1/XA4/MP2/a_216_n18# 0.01fF
C3585 XDAC2/XC1/XRES1B/B XDAC2/XC64a<0>/XRES16/B 0.05fF
C3586 XA4/XA3/MP1/a_216_n18# AVDD 0.07fF
C3587 XDAC1/XC1/XRES8/B XB1/XA4/GNG 0.33fF
C3588 XDAC1/XC1/XRES16/B XB1/XA3/B 0.17fF
C3589 XA20/XA9/A XA20/XA10/MN1/a_324_n18# 0.01fF
C3590 XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C3591 XA7/EN AVDD 4.92fF
C3592 XA5/XA9/Y XA5/XA11/MP0/a_216_n18# 0.08fF
C3593 XA8/XA12/A AVSS 0.42fF
C3594 XA8/XA1/XA4/MP2/S XA8/XA4/A 0.05fF
C3595 XA7/XA1/XA1/MP0/a_216_n18# XA7/EN 0.01fF
C3596 XA4/XA1/XA4/MP1/S XA20/CPO 0.02fF
C3597 XA1/XA2/MP1/a_216_n18# VREF 0.02fF
C3598 XA7/XA9/A XA7/XA9/MN1/a_324_n18# 0.07fF
C3599 XA5/CEO AVDD 0.71fF
C3600 XA1/EN XA0/XA1/XA4/MN0/a_324_n18# 0.07fF
C3601 XA4/XA2/MN0/a_324_n18# XA4/EN 0.07fF
C3602 XA3/XA1/XA1/MP0/a_216_n18# XA3/EN 0.01fF
C3603 D<1> XA3/CN1 0.04fF
C3604 XA4/EN XA20/CNO 1.01fF
C3605 XA5/XA4/MP1/a_216_n18# XA5/XA4/MP2/a_216_n18# 0.01fF
C3606 XA5/XA4/MN0/a_324_n18# AVSS 0.01fF
C3607 XB1/CKN XB1/XA3/MP0/a_216_n18# 0.08fF
C3608 XA0/XA11/A AVDD 0.45fF
C3609 XA5/XA11/A XA5/XA11/MP0/a_216_n18# 0.07fF
C3610 XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MP2/a_216_n18# 0.01fF
C3611 XA6/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C3612 D<2> D<1> 3.28fF
C3613 XA4/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C3614 XA1/EN AVSS 1.13fF
C3615 XA7/XA6/MN1/S AVSS 0.15fF
C3616 XA4/XA5/MP3/a_216_n18# AVDD 0.07fF
C3617 XA4/XA5/MN3/a_324_n18# XA4/CP0 0.15fF
C3618 XA6/XA2/A XA6/CN1 0.57fF
C3619 XA0/CEO XA0/XA13/MP1/a_216_n18# 0.01fF
C3620 XDAC1/XC1/XRES2/B SARP 3.05fF
C3621 XA5/XA1/XA5/MN1/S EN 0.01fF
C3622 SAR_IN XB2/M1/a_324_n18# 0.01fF
C3623 XA2/CN0 XA20/CNO 0.05fF
C3624 XA6/CN0 XA2/CN1 0.45fF
C3625 D<1> XA7/CN0 2.67fF
C3626 XA1/XA4/A XA1/CN0 0.10fF
C3627 XA8/XA2/MP1/a_216_n18# AVDD 0.08fF
C3628 XA2/EN XA1/XA1/XA1/MP3/a_216_n18# 0.01fF
C3629 XA7/XA3/MP1/a_216_n18# AVDD 0.07fF
C3630 XA20/XA9/Y XA20/XA3/MP0/a_216_n18# 0.07fF
C3631 XA4/XA5/MP1/a_216_n18# XA4/CN0 0.02fF
C3632 XB2/XA3/B XB2/XCAPB1/XCAPB2/m3_9828_132# 0.21fF
C3633 XB2/XA1/Y XB2/XA2/MP0/G 0.01fF
C3634 D<1> D<3> 1.30fF
C3635 XA7/CEO XA8/XA12/MN0/a_324_n18# 0.07fF
C3636 XA6/XA6/MP0/a_216_n18# XA6/CP0 0.08fF
C3637 XA1/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C3638 XA4/XA9/Y VREF 0.03fF
C3639 XA0/CP0 XA1/CN0 0.01fF
C3640 XA5/EN XA5/XA2/MN0/a_324_n18# 0.07fF
C3641 XA20/XA3/MP5/a_216_n18# XA20/XA3/MP4/a_216_n18# 0.01fF
C3642 XA1/XA11/MP1/S VREF 0.01fF
C3643 XA0/XA1/XA1/MP0/a_216_n18# XA0/XA1/XA1/MP1/a_216_n18# 0.01fF
C3644 XA3/XA1/XA4/MN1/S XA4/EN 0.01fF
C3645 XB1/XCAPB1/XCAPB1/m3_324_308# XB1/XA3/B 0.02fF
C3646 XA3/EN XA2/XA1/XA4/MP1/S 0.02fF
C3647 XA4/XA9/MP1/a_216_334# AVDD 0.09fF
C3648 XA20/CNO SARN 0.03fF
C3649 XA8/XA1/XA2/MN0/a_324_n18# XA8/XA1/XA4/MN0/a_324_n18# 0.01fF
C3650 XA3/XA3/MP3/a_216_n18# XA3/XA3/MP2/a_216_n18# 0.01fF
C3651 XA2/XA6/MP3/S VREF 0.02fF
C3652 XA8/XA5/MP2/a_216_n18# XA8/CP0 0.15fF
C3653 D<1> XA7/XA1/XA1/MN2/S 0.01fF
C3654 XA2/XA1/XA2/Y XA2/XA1/XA5/MN0/a_324_n18# 0.02fF
C3655 XDAC2/X16ab/XRES1A/B XDAC2/X16ab/XRES4/B 0.29fF
C3656 XDAC2/X16ab/XRES2/B XDAC2/X16ab/XRES1B/B 0.23fF
C3657 XA0/DONE AVSS 0.15fF
C3658 XDAC2/XC128a<1>/XRES2/B AVSS 3.71fF
C3659 SARP XB1/M6/a_324_n18# 0.02fF
C3660 XDAC1/X16ab/XRES2/B AVSS 3.71fF
C3661 XA7/XA12/MN0/a_324_n18# XA7/XA13/MN1/a_324_n18# 0.01fF
C3662 XDAC1/XC64b<1>/XRES8/B AVSS 9.08fF
C3663 D<2> XA3/CN1 0.03fF
C3664 XA5/XA1/XA2/Y AVSS 0.31fF
C3665 XA7/XA4/MN3/a_324_n18# XA7/XA4/A 0.15fF
C3666 XA6/XA1/XA4/MN1/S AVSS 0.10fF
C3667 XA4/XA9/B AVDD 0.79fF
C3668 XA3/CN0 D<5> 0.50fF
C3669 XDAC2/XC128a<1>/XRES2/B XDAC2/XC128a<1>/XRES1B/B 0.23fF
C3670 XA1/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C3671 XA8/CN1 XA20/XA3/CO 0.05fF
C3672 XDAC1/X16ab/XRES2/B XDAC1/X16ab/XRES1B/B 0.23fF
C3673 XA7/CN0 XA3/CN1 0.05fF
C3674 XB1/XCAPB1/XCAPB3/m3_252_308# XB1/XA4/GNG 0.13fF
C3675 XA2/CN1 XA2/XA3/MN3/a_324_n18# 0.15fF
C3676 XA1/EN CK_SAMPLE 0.09fF
C3677 XA8/XA3/MP3/a_216_n18# AVDD 0.07fF
C3678 XA7/XA6/MN1/S CK_SAMPLE 0.05fF
C3679 XA1/XA1/XA5/MN1/a_324_n18# XA20/CNO 0.07fF
C3680 XA7/XA13/MP1/a_216_n18# AVDD 0.13fF
C3681 XA20/XA2/MP5/a_216_n18# XA20/XA3/CO 0.15fF
C3682 XDAC1/XC32a<0>/XRES8/B AVSS 9.20fF
C3683 XA4/CN0 AVDD 5.33fF
C3684 XDAC1/XC64b<1>/XRES4/B XDAC1/X16ab/XRES4/B 0.10fF
C3685 XDAC1/XC64b<1>/XRES8/B XDAC1/X16ab/XRES1B/B 0.02fF
C3686 XA7/EN XA6/XA1/XA1/MP3/a_216_n18# 0.02fF
C3687 XB2/XA3/MP2/a_216_n18# XB2/XA3/MP0/a_216_334# 0.01fF
C3688 EN XA2/XA1/XA5/MP2/S 0.04fF
C3689 XA8/XA9/MP0/a_216_n18# XA8/XA9/MP1/a_216_n18# 0.01fF
C3690 XA8/XA4/MP1/a_216_n18# AVDD 0.07fF
C3691 XA0/XA11/MN1/a_324_n18# XA0/XA12/A 0.01fF
C3692 XB1/XA5/MN1/a_324_n18# XB1/XA2/MP0/G 0.06fF
C3693 XA2/XA2/A AVSS 0.23fF
C3694 XA8/XA12/MP0/a_216_n18# XA8/XA12/A 0.07fF
C3695 XA0/XA4/A XA0/XA4/MN1/a_324_n18# 0.15fF
C3696 XA3/XA1/XA5/MN1/S AVSS 0.12fF
C3697 XA0/XA12/MN0/a_324_n18# XA0/CEIN 0.07fF
C3698 D<3> XA3/CN1 0.03fF
C3699 XA7/XA1/XA4/MP1/S XA7/XA1/XA4/MN1/S 0.01fF
C3700 XA5/CN0 AVDD 4.40fF
C3701 D<2> XA7/CN0 0.17fF
C3702 XB2/XA4/GNG XB2/XA4/MP1/a_216_334# 0.02fF
C3703 EN XA1/EN 1.06fF
C3704 XB2/XA3/B XDAC2/XC1/XRES16/B 0.17fF
C3705 XA0/XA1/XA0/MP1/a_216_n18# AVDD 0.15fF
C3706 XA0/XA1/XA5/MN1/a_324_n18# XA0/XA1/XA2/Y 0.09fF
C3707 XA1/XA1/XA1/MP3/S XA2/EN 0.10fF
C3708 XA4/XA6/MP0/a_216_n18# VREF 0.01fF
C3709 XA5/XA1/XA1/MP1/a_216_n18# AVDD 0.08fF
C3710 XA0/XA9/Y XA0/XA12/A 0.02fF
C3711 XA3/CP0 XA2/CN1 0.03fF
C3712 XB2/XA1/Y XB2/XA4/MN1/a_324_334# 0.08fF
C3713 D<1> XA8/EN 0.47fF
C3714 XA4/XA9/B XA4/XA9/MN1/S 0.02fF
C3715 XA3/XA3/MP2/a_216_n18# AVDD 0.07fF
C3716 XA6/XA4/MP2/a_216_n18# AVDD 0.07fF
C3717 XA7/XA1/XA1/MP3/G XA20/CPO 0.15fF
C3718 XA4/CN0 XA4/XA1/XA2/Y 0.02fF
C3719 XDAC2/XC1/XRES16/B AVSS 15.88fF
C3720 XA6/XA13/MP1/a_216_n18# AVDD 0.13fF
C3721 XDAC1/XC32a<0>/XRES16/B XDAC1/XC64a<0>/XRES8/B 0.03fF
C3722 XA7/XA9/B XA7/XA6/MP1/S 0.07fF
C3723 XB2/XCAPB1/XCAPB3/m3_324_308# XB2/XA3/B 0.02fF
C3724 D<2> D<3> 2.96fF
C3725 XA0/XA3/MN1/a_324_n18# XA0/XA3/MN2/a_324_n18# 0.01fF
C3726 XA5/CP0 XA5/XA4/MN1/a_324_n18# 0.03fF
C3727 XA1/XA5/MP0/a_216_n18# VREF 0.02fF
C3728 XA8/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C3729 XA8/XA4/MP3/a_216_n18# XA8/XA4/A 0.15fF
C3730 XA6/XA4/A XA20/CNO 0.18fF
C3731 XDAC1/XC0/XRES16/B SARP 21.65fF
C3732 XA7/XA4/MP3/a_216_n18# VREF 0.03fF
C3733 XA7/CN0 D<3> 0.15fF
C3734 XA7/XA9/A XA7/XA9/Y 0.04fF
C3735 XA0/CN0 XA1/CN1 1.21fF
C3736 DONE AVDD 2.20fF
C3737 XA7/XA3/MP3/a_216_n18# XA7/CN1 0.15fF
C3738 XA6/XA9/B XA6/XA9/MN1/a_324_334# 0.07fF
C3739 XA2/XA9/Y XA2/XA9/MP1/a_216_334# 0.07fF
C3740 XB2/XA1/Y XB2/CKN 0.08fF
C3741 XA5/XA11/MP1/a_216_n18# XA4/CEO 0.07fF
C3742 XDAC1/XC0/XRES1A/B AVSS 2.94fF
C3743 XA3/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C3744 XA7/XA8/MP0/a_216_n18# XA7/XA9/A 0.07fF
C3745 XA4/XA1/XA5/MP1/S VREF 0.02fF
C3746 XDAC1/XC128b<2>/XRES1B/B SARP 1.79fF
C3747 XA5/XA6/MP3/a_216_n18# AVDD 0.08fF
C3748 XA0/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C3749 XA6/EN XA5/XA1/XA5/MP2/S 0.02fF
C3750 VREF XA3/XA4/A 0.37fF
C3751 XA5/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C3752 XA20/XA1/MP0/S XA20/XA1/MN2/a_324_n18# 0.01fF
C3753 XDAC2/XC0/XRES4/B SARN 6.39fF
C3754 XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C3755 D<0> XA20/XA3a/A 0.03fF
C3756 XDAC2/XC128a<1>/XRES1A/B XDAC2/XC32a<0>/XRES4/B 0.01fF
C3757 VREF XA0/CEO 0.26fF
C3758 XA5/XA7/MP0/a_216_n18# AVDD 0.09fF
C3759 XA4/XA1/XA5/MN2/a_324_n18# XA4/EN 0.08fF
C3760 XA2/CN0 XA2/XA1/XA2/Y 0.02fF
C3761 XA6/EN XA5/XA6/MP3/S 0.02fF
C3762 XA6/CN0 VREF 0.69fF
C3763 XA5/XA1/XA2/Y EN 0.07fF
C3764 XA7/EN XA7/XA2/A 0.09fF
C3765 XDAC2/XC1/XRES2/B XDAC2/XC64a<0>/XRES2/B 0.05fF
C3766 XA7/XA2/MP1/a_216_n18# AVDD 0.08fF
C3767 XA3/XA1/XA5/MP2/S EN 0.04fF
C3768 XA20/XA9/Y XA20/CNO 0.07fF
C3769 XA2/XA5/MP2/a_216_n18# AVDD 0.07fF
C3770 XA1/XA4/MP3/a_216_n18# VREF 0.03fF
C3771 XA2/EN XA1/XA1/XA4/MN1/S 0.01fF
C3772 XA0/XA13/MN1/a_324_334# XA0/XA13/MN1/a_324_n18# 0.01fF
C3773 XA4/XA2/A XA4/XA3/MN0/a_324_n18# 0.07fF
C3774 XA1/XA11/MP0/a_216_n18# XA1/XA11/MP1/a_216_n18# 0.01fF
C3775 XA6/XA11/MP0/a_216_n18# XA6/XA9/MP1/a_216_334# 0.01fF
C3776 XA6/CP0 AVDD 1.31fF
C3777 XB1/M7/a_324_n18# XB1/M6/a_324_n18# 0.01fF
C3778 D<7> XA3/CP0 0.05fF
C3779 XA5/CP0 XA4/CP0 0.03fF
C3780 XDAC1/XC1/XRES1A/B XB1/XA3/B 0.21fF
C3781 XA20/XA3/MN0/a_324_n18# XA20/XA3a/MN3/a_324_n18# 0.01fF
C3782 XA3/XA6/MN0/a_324_n18# AVSS 0.01fF
C3783 XA4/XA1/XA2/Y XA4/XA1/XA4/MN0/a_324_n18# 0.02fF
C3784 XA2/XA2/A EN 0.13fF
C3785 XDAC1/XC32a<0>/XRES2/B XDAC1/XC128a<1>/XRES2/B 0.05fF
C3786 XA3/XA8/MP0/a_216_n18# XA3/XA9/MP0/a_216_n18# 0.01fF
C3787 XA3/XA9/B XA3/XA9/MN0/a_324_n18# 0.01fF
C3788 XA1/XA8/MP0/a_216_n18# XA1/XA9/MP0/a_216_n18# 0.01fF
C3789 XA3/XA1/XA5/MN1/S EN 0.01fF
C3790 XA3/XA1/XA5/MP0/a_216_n18# EN 0.16fF
C3791 XDAC2/XC128b<2>/XRES16/B AVSS 16.02fF
C3792 XA4/XA9/MP0/a_216_n18# XA4/XA9/A 0.14fF
C3793 D<2> XA8/EN 0.02fF
C3794 XA7/XA12/A XA7/XA11/MP1/S 0.06fF
C3795 XDAC2/XC64b<1>/XRES4/B AVSS 5.49fF
C3796 XDAC2/XC1/XRES4/B XDAC2/XC64a<0>/XRES4/B 0.10fF
C3797 XA8/XA4/MN0/a_324_n18# XA8/XA4/MN1/a_324_n18# 0.01fF
C3798 XA3/XA1/XA5/MP1/S EN 0.03fF
C3799 XA4/XA9/B XA5/EN 0.07fF
C3800 XA4/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C3801 XA5/XA1/XA4/MN1/S AVSS 0.10fF
C3802 XDAC1/XC128a<1>/XRES8/B SARP 11.94fF
C3803 XA4/XA4/A XA4/XA3/MN3/a_324_n18# 0.01fF
C3804 XA2/XA1/XA2/Y XA2/XA1/XA4/MN1/S 0.05fF
C3805 XA8/XA12/MN0/a_324_n18# AVSS 0.01fF
C3806 XA3/XA12/A XA3/XA12/MN0/a_324_n18# 0.09fF
C3807 XA8/EN XA7/CN0 0.20fF
C3808 XA0/XA9/A XA0/XA9/B 0.29fF
C3809 XA6/XA11/MP0/a_216_n18# AVDD 0.09fF
C3810 XDAC2/XC128b<2>/XRES4/B SARN 6.32fF
C3811 XDAC2/XC128a<1>/XRES16/B AVSS 16.02fF
C3812 XDAC2/XC128b<2>/XRES16/B XDAC2/XC128a<1>/XRES1B/B 0.05fF
C3813 XA1/XA1/XA4/MP2/S EN 0.03fF
C3814 XA4/CN0 XA5/EN 0.15fF
C3815 XA20/XA9/A XA20/CNO 0.07fF
C3816 XA0/XA11/MP0/a_216_n18# AVDD 0.09fF
C3817 XA2/XA4/A XA2/XA1/XA4/MN2/S 0.06fF
C3818 XDAC1/XC64a<0>/XRES2/B AVSS 3.71fF
C3819 XA0/XA4/MP3/a_216_n18# AVDD 0.07fF
C3820 XB1/XA4/GNG XB1/XA4/MP1/a_216_334# 0.02fF
C3821 XA20/CPO XA0/XA1/XA1/MN3/a_324_n18# 0.08fF
C3822 XA7/XA4/MP2/a_216_n18# VREF 0.03fF
C3823 XA1/XA11/A AVDD 0.45fF
C3824 XDAC2/XC128a<1>/XRES1B/B XDAC2/XC128a<1>/XRES16/B 0.12fF
C3825 XA1/XA9/MN1/a_324_334# XA1/XA9/MN1/a_324_n18# 0.01fF
C3826 XA2/XA11/A XA2/XA11/MP1/a_216_n18# 0.08fF
C3827 XA8/XA11/MP0/a_216_n18# XA8/XA9/Y 0.08fF
C3828 XA5/CN0 XA5/EN 0.11fF
C3829 XA7/XA1/XA1/MP3/G XA7/XA1/XA2/MN0/a_324_n18# 0.06fF
C3830 XA3/XA1/XA2/Y AVSS 0.27fF
C3831 XA20/XA1/MP0/S SARN 0.03fF
C3832 XA0/XA2/A XA0/XA2/MN0/a_324_n18# 0.08fF
C3833 XA0/XA1/XA5/MP2/S VREF 0.03fF
C3834 XA3/XA9/A XA3/XA9/MN1/a_324_n18# 0.07fF
C3835 XA6/XA3/MP3/a_216_n18# XA6/CN1 0.15fF
C3836 XA2/XA2/A XA2/XA2/MP1/a_216_n18# 0.15fF
C3837 XA0/XA12/A XA0/CEIN 0.13fF
C3838 XA5/XA12/A XA5/XA11/MP1/S 0.06fF
C3839 XA7/XA4/MP0/a_216_n18# AVDD 0.08fF
C3840 XA4/XA2/A XA4/XA2/MN2/a_324_n18# 0.15fF
C3841 EN XA0/XA1/XA5/MP1/a_216_n18# 0.16fF
C3842 XA20/XA11/MN1/a_324_n18# XA20/XA11/Y 0.02fF
C3843 XA8/XA2/MN0/a_324_n18# XA8/XA2/A 0.08fF
C3844 XB2/XA7/MP1/a_216_n18# XB2/XA1/MP0/G 0.08fF
C3845 D<5> XA20/CNO 0.06fF
C3846 XA2/XA11/A XA2/XA11/MN1/a_324_n18# 0.07fF
C3847 XA0/XA1/XA4/MN2/S AVSS 0.06fF
C3848 XA1/XA6/MP0/a_216_n18# VREF 0.01fF
C3849 XA3/EN XA2/XA1/XA1/MP3/a_216_n18# 0.02fF
C3850 XB1/XA4/MP1/a_216_n18# XB1/XA4/GNG 0.02fF
C3851 XA8/EN XA7/XA1/XA1/MN2/S 0.11fF
C3852 XDAC1/XC0/XRES1A/B XDAC1/XC0/XRES2/B 0.25fF
C3853 SAR_IP XB1/M4/a_324_n18# 0.02fF
C3854 AVDD XA8/XA6/MN1/S 0.01fF
C3855 XB2/XA3/MN2/a_324_n18# XB2/XA3/B 0.01fF
C3856 XA2/XA1/XA4/MP1/S XA2/XA1/XA4/MP2/S 0.04fF
C3857 XA3/XA2/MN1/a_324_n18# XA3/CN1 0.03fF
C3858 D<6> XA1/CN1 0.05fF
C3859 XA1/XA4/A XA1/XA5/MN0/a_324_n18# 0.07fF
C3860 XA2/EN XA20/CPO 0.76fF
C3861 XA5/XA9/MN1/S AVDD 0.01fF
C3862 XB2/XA1/Y XA0/CEIN 0.07fF
C3863 XA7/XA1/XA4/MP1/S XA20/CPO 0.03fF
C3864 XA1/XA9/B XA1/XA6/MN3/S 0.09fF
C3865 XA5/XA12/A XA5/XA12/MN0/a_324_n18# 0.09fF
C3866 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MP2/S 0.04fF
C3867 XA3/CP0 VREF 0.83fF
C3868 XA20/XA11/MP1/a_216_n18# XA20/XA12/MP0/a_216_n18# 0.01fF
C3869 XA8/ENO XA20/XA2/N2 0.01fF
C3870 XB2/XA7/MP1/a_216_334# XB2/XA7/MP1/a_216_n18# 0.01fF
C3871 XA4/XA11/MN0/a_324_n18# AVSS 0.01fF
C3872 XA3/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C3873 XA20/CNO XA3/XA1/XA1/MN2/S 0.03fF
C3874 XA20/XA3a/MN2/a_324_n18# XA20/XA3a/MN1/a_324_n18# 0.01fF
C3875 XA2/EN XA1/XA7/MP0/a_216_n18# 0.07fF
C3876 XA6/EN XA5/XA1/XA4/MN2/S 0.01fF
C3877 XB2/XA3/MN0/a_324_n18# AVSS 0.01fF
C3878 XA1/XA6/MP3/a_216_n18# XA1/XA7/MP0/a_216_n18# 0.01fF
C3879 XA1/CEO XA1/XA9/Y 0.03fF
C3880 AVDD XA20/XA2/MP6/a_216_334# 0.09fF
C3881 XDAC1/X16ab/XRES1A/B XDAC1/X16ab/XRES2/B 0.25fF
C3882 D<3> XA5/XA3/MP2/a_216_n18# 0.01fF
C3883 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MP3/a_216_n18# 0.07fF
C3884 XA5/EN XA4/XA1/XA4/MN0/a_324_n18# 0.07fF
C3885 SARP XB1/XA1/Y 0.02fF
C3886 XA2/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C3887 XA3/XA2/A XA3/XA4/A 0.14fF
C3888 XA3/XA1/XA5/MN2/S XA20/CNO 0.01fF
C3889 XDAC2/X16ab/XRES1B/B XDAC2/X16ab/XRES16/B 0.12fF
C3890 EN XA2/XA1/XA1/MP1/a_216_n18# 0.08fF
C3891 XA2/XA3/MP3/a_216_n18# XA2/XA4/MP0/a_216_n18# 0.01fF
C3892 XA8/ENO XA20/XA3a/A 0.15fF
C3893 VREF XA3/XA4/MP1/a_216_n18# 0.02fF
C3894 XA0/XA9/B AVDD 0.79fF
C3895 D<1> XA7/XA6/MP3/S 0.02fF
C3896 XA7/XA4/A AVSS 1.11fF
C3897 XA1/XA1/XA2/Y XA1/XA1/XA4/MP1/S 0.01fF
C3898 SARP XB1/CKN 0.05fF
C3899 XA3/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C3900 D<1> XA7/XA7/MP0/a_216_n18# 0.08fF
C3901 XA1/XA2/A XA1/XA2/MN1/a_324_n18# 0.15fF
C3902 XA3/CN0 AVDD 4.37fF
C3903 XA7/XA1/XA5/MP1/S AVDD 0.13fF
C3904 XA4/CN0 XDAC2/XC32a<0>/XRES16/B 0.02fF
C3905 XB1/XA4/MN1/a_324_334# XB1/XA1/Y 0.08fF
C3906 XA7/XA6/MP1/S CK_SAMPLE 0.03fF
C3907 XA6/XA11/MP1/a_216_n18# XA6/XA11/A 0.08fF
C3908 XB1/M4/G XB1/XA4/GNG 0.25fF
C3909 XA1/CN1 SARP 0.20fF
C3910 XB1/XA1/MP0/G XB1/XA7/MP1/a_216_n18# 0.08fF
C3911 XA4/XA1/XA4/MN1/a_324_n18# XA4/XA1/XA4/MN2/a_324_n18# 0.01fF
C3912 XA6/XA11/MN0/a_324_n18# XA6/XA11/A 0.09fF
C3913 XDAC2/XC64b<1>/XRES1A/B XDAC2/X16ab/XRES8/B 0.03fF
C3914 D<1> XA7/CN1 0.43fF
C3915 XA6/EN XA6/XA1/XA1/MN2/S 0.05fF
C3916 XA8/XA3/MP1/a_216_n18# XA8/CN1 0.15fF
C3917 EN XA0/XA1/XA1/MP1/a_216_n18# 0.08fF
C3918 XA1/XA12/A AVSS 0.39fF
C3919 XA3/XA1/XA4/MN2/S AVSS 0.06fF
C3920 XA2/XA11/MN1/a_324_n18# AVSS 0.01fF
C3921 XA3/XA1/XA4/MP1/S XA3/XA1/XA4/MN1/S 0.01fF
C3922 D<0> XA8/XA3/MN3/a_324_n18# 0.02fF
C3923 AVDD XA20/XA3/MP0/a_216_n18# 0.09fF
C3924 XA4/XA1/XA5/MP2/S VREF 0.03fF
C3925 XA3/XA4/MP0/a_216_n18# XA3/XA4/A 0.07fF
C3926 XA5/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C3927 XA5/XA2/A AVSS 0.28fF
C3928 XA5/CN0 XDAC2/XC32a<0>/XRES16/B 0.02fF
C3929 XA5/XA6/MN0/a_324_n18# AVSS 0.01fF
C3930 XA6/XA5/MP0/a_216_n18# XA6/CP0 0.07fF
C3931 XA7/XA4/MP1/a_216_n18# VREF 0.02fF
C3932 XA4/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C3933 EN XA3/XA1/XA2/Y 0.07fF
C3934 XA0/XA1/XA1/MP3/S XA0/XA1/XA1/MP2/S 0.04fF
C3935 CK_SAMPLE_BSSW XB1/XA3/B 0.05fF
C3936 XA5/XA4/A XA5/XA1/XA5/MN1/S 0.02fF
C3937 EN XA2/XA1/XA4/MP2/a_216_n18# 0.15fF
C3938 XA0/XA7/MN0/a_324_n18# AVSS 0.01fF
C3939 XA1/XA9/B XA1/XA8/MN0/a_324_n18# 0.01fF
C3940 D<0> XA8/XA6/MP1/a_216_n18# 0.01fF
C3941 SARN XB1/M8/a_324_n18# 0.02fF
C3942 XA6/XA2/A XA6/XA2/MP0/a_216_n18# 0.08fF
C3943 AVDD XB1/XA4/GNG 4.07fF
C3944 EN XA0/XA1/XA4/MN2/S 0.02fF
C3945 XA8/XA4/MP0/a_216_n18# XA8/CN1 0.08fF
C3946 D<7> XA1/XA6/MP1/a_216_n18# 0.01fF
C3947 XA20/XA13/MP1/a_216_n18# AVDD 0.13fF
C3948 XA20/XA2/MP0/a_216_n18# XA20/XA9/Y 0.07fF
C3949 XA4/XA2/MN1/a_324_n18# XA4/XA2/MN0/a_324_n18# 0.01fF
C3950 XA20/XA3a/A XA8/CN0 0.02fF
C3951 XA2/CN1 XA1/EN 0.08fF
C3952 XB2/XA3/B XB2/XCAPB1/XCAPB2/m3_252_308# 0.02fF
C3953 XDAC2/XC64b<1>/XRES4/B XDAC2/XC0/XRES1A/B 0.01fF
C3954 XDAC2/XC64b<1>/XRES4/B XDAC2/XC64b<1>/XRES8/B 2.60fF
C3955 XA6/EN XA5/XA1/XA4/MP2/S 0.02fF
C3956 XA4/XA6/MN2/a_324_n18# AVSS 0.01fF
C3957 XA1/XA4/MP0/a_216_n18# XA1/CN1 0.08fF
C3958 XDAC1/XC32a<0>/XRES16/B XDAC1/XC64a<0>/XRES1B/B 0.05fF
C3959 XA0/CN0 AVSS 2.03fF
C3960 XDAC1/XC128b<2>/XRES4/B SARP 6.32fF
C3961 XA7/XA5/MP2/a_216_n18# VREF 0.03fF
C3962 AVDD XA20/XA4/MP2_DMY/a_216_n18# 0.24fF
C3963 XA20/XA2a/MP2/a_216_n18# XA20/XA3/CO 0.16fF
C3964 XA4/XA2/A XA3/XA4/A 0.03fF
C3965 XA20/XA12/Y XA20/XA11/MP1/S 0.04fF
C3966 XA1/XA11/A XA1/XA11/MN1/a_324_n18# 0.07fF
C3967 D<6> XA2/XA4/MP0/a_216_n18# 0.01fF
C3968 XA7/XA2/MP1/a_216_n18# XA7/XA2/A 0.15fF
C3969 XA1/XA11/A XA1/XA9/A 0.01fF
C3970 XA4/XA1/XA5/MN2/S XA4/XA4/A 0.02fF
C3971 XDAC1/XC64b<1>/XRES16/B XDAC1/X16ab/XRES16/B 0.41fF
C3972 XDAC2/XC128b<2>/XRES1B/B XDAC2/XC128b<2>/XRES4/B 1.64fF
C3973 XDAC2/XC128b<2>/XRES2/B XDAC2/XC128b<2>/XRES8/B 1.58fF
C3974 XDAC2/XC0/XRES2/B XDAC2/XC0/XRES4/B 0.55fF
C3975 XA8/XA3/MN2/a_324_n18# XA8/XA3/MN3/a_324_n18# 0.01fF
C3976 XA5/CP0 AVDD 1.31fF
C3977 XA5/XA6/MP1/a_216_n18# AVDD 0.08fF
C3978 XA3/XA2/MP1/a_216_n18# XA3/XA2/MP0/a_216_n18# 0.01fF
C3979 XA1/XA12/MN0/a_324_n18# XA0/CEO 0.07fF
C3980 XDAC1/XC64b<1>/XRES2/B XDAC1/XC64b<1>/XRES1A/B 0.25fF
C3981 XB2/XA3/MN0/a_324_n18# XB2/XA0/MN0/a_324_n18# 0.01fF
C3982 XB1/XCAPB1/XCAPB3/m3_9756_132# XB1/XA3/B 0.07fF
C3983 XA5/CP0 XA5/XA4/MN2/a_324_n18# 0.01fF
C3984 XA8/XA13/MN1/a_324_334# AVSS 0.10fF
C3985 XA0/XA8/MN0/a_324_n18# XA0/XA9/B 0.01fF
C3986 XA2/XA9/Y XA2/XA11/MN0/a_324_n18# 0.07fF
C3987 XA1/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C3988 D<2> XA7/CN1 0.01fF
C3989 XA7/XA1/XA5/MN1/S AVDD 0.02fF
C3990 EN XA5/XA1/XA4/MP1/S 0.02fF
C3991 XA8/XA12/A XA8/XA9/B 0.01fF
C3992 XA7/XA4/A EN 0.09fF
C3993 XA20/XA3a/A XA20/XA3a/MP1/a_216_n18# 0.16fF
C3994 XB2/M3/a_324_n18# SARN 0.01fF
C3995 XA5/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C3996 XA0/XA11/MP1/a_216_n18# XA0/XA12/MP0/a_216_n18# 0.01fF
C3997 XA4/XA11/MP0/a_216_n18# AVDD 0.09fF
C3998 XA3/XA2/A XA3/CP0 0.04fF
C3999 XA20/XA1/MP0/S XA20/XA9/A 0.13fF
C4000 EN XA2/XA1/XA5/MP1/a_216_n18# 0.16fF
C4001 XA5/XA6/MP0/a_216_n18# XA5/XA5/MP3/a_216_n18# 0.01fF
C4002 XA7/CN0 XA7/CN1 0.08fF
C4003 XA20/XA3/MN6/a_324_n18# XA20/XA3a/A 0.08fF
C4004 XA1/XA2/MP0/a_216_n18# XA1/XA2/A 0.08fF
C4005 XA2/EN XA1/CP0 0.16fF
C4006 XA8/XA1/XA1/MP3/S AVSS 0.03fF
C4007 VREF XA20/XA3/CO 0.32fF
C4008 XA5/XA4/MN0/a_324_n18# XA5/XA4/A 0.09fF
C4009 D<4> D<8> 0.10fF
C4010 XA0/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C4011 XA1/XA6/MN0/a_324_n18# XA1/XA5/MN3/a_324_n18# 0.01fF
C4012 XA7/XA1/XA4/MP2/S AVDD 0.11fF
C4013 XA3/XA2/MN0/a_324_n18# XA3/XA2/MN1/a_324_n18# 0.01fF
C4014 XA5/XA2/A EN 0.12fF
C4015 XA4/XA9/B XA3/XA9/B 0.07fF
C4016 XA5/XA2/A XA5/XA3/MN0/a_324_n18# 0.07fF
C4017 XA5/XA1/XA5/MN0/a_324_n18# XA5/XA1/XA2/Y 0.02fF
C4018 XA20/CPO XA2/XA1/XA1/MN3/a_324_n18# 0.08fF
C4019 D<1> XA0/CP0 0.05fF
C4020 XDAC1/XC1/XRES1B/B AVSS 2.94fF
C4021 XA6/XA12/MN0/a_324_n18# AVSS 0.01fF
C4022 XA6/XA1/XA4/MP1/a_216_n18# XA6/XA1/XA4/MP0/a_216_n18# 0.01fF
C4023 XA4/XA6/MN0/a_324_n18# AVSS 0.01fF
C4024 XA0/XA12/A XA0/XA12/MN0/a_324_n18# 0.09fF
C4025 XA7/XA6/MP0/a_216_n18# XA7/CP0 0.08fF
C4026 XA1/XA13/MN1/a_324_334# AVSS 0.10fF
C4027 XA2/XA7/MN0/a_324_n18# XA3/EN 0.08fF
C4028 D<7> XA1/EN 0.09fF
C4029 XA3/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C4030 XA5/CN1 AVSS 0.80fF
C4031 XA4/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C4032 XA8/XA1/XA4/MP1/S XA8/XA1/XA4/MP2/S 0.04fF
C4033 XDAC1/XC1/XRES2/B XB1/XA4/GNG 0.19fF
C4034 XA20/XA2/MN6/a_324_n18# XA20/XA2/MN5/a_324_n18# 0.01fF
C4035 XA0/CN0 CK_SAMPLE 0.09fF
C4036 XA2/XA2/A XA2/CN1 0.62fF
C4037 XA7/CN0 XA7/XA5/MP1/a_216_n18# 0.02fF
C4038 XA7/XA2/MN0/a_324_n18# XA7/XA2/A 0.08fF
C4039 XA6/XA1/XA4/MN2/S XA6/XA1/XA2/Y 0.05fF
C4040 XA1/XA2/MN1/a_324_n18# XA1/CN1 0.03fF
C4041 XA2/XA1/XA5/MP1/S XA2/XA1/XA5/MN1/S 0.01fF
C4042 XA8/XA4/MP2/a_216_n18# XA8/XA4/MP1/a_216_n18# 0.01fF
C4043 XA2/DONE AVSS 0.15fF
C4044 XA2/XA12/A XA2/XA11/MN1/a_324_n18# 0.01fF
C4045 XA2/XA2/MP3/a_216_n18# XA2/XA2/MP2/a_216_n18# 0.01fF
C4046 XA1/XA1/XA1/MP2/a_216_n18# XA1/XA1/XA1/MP3/G 0.01fF
C4047 XA1/XA6/MP1/S AVDD 0.12fF
C4048 XA2/CP0 D<8> 0.03fF
C4049 XA2/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C4050 XDAC2/X16ab/XRES2/B AVSS 3.71fF
C4051 XA20/XA4/MP2_DMY/a_216_n18# XA20/XA4/MP3_DMY/a_216_n18# 0.01fF
C4052 XA4/DONE AVSS 0.15fF
C4053 XA2/CP0 XA2/XA5/MP1/a_216_n18# 0.15fF
C4054 XA4/XA3/MP0/a_216_n18# XA4/CN1 0.07fF
C4055 EN XA0/CN0 0.08fF
C4056 SARN XDAC2/XC32a<0>/XRES1B/B 1.79fF
C4057 XA3/XA4/MP0/a_216_n18# XA3/XA4/MP1/a_216_n18# 0.01fF
C4058 XA5/XA3/MP3/a_216_n18# VREF 0.03fF
C4059 XA8/XA3/MP0/a_216_n18# AVDD 0.08fF
C4060 XA7/XA4/A XA8/CN1 0.04fF
C4061 XA8/XA4/MN1/a_324_n18# XA8/XA4/A 0.15fF
C4062 XA2/CP0 XA2/XA4/A 0.57fF
C4063 XA1/XA1/XA4/MN2/S XA1/XA4/A 0.06fF
C4064 XA20/CNO AVDD 8.74fF
C4065 XDAC1/XC128b<2>/XRES1B/B XDAC1/X16ab/XRES8/B 0.02fF
C4066 XA8/XA1/XA5/MP2/S XA8/XA1/XA5/MN2/S 0.01fF
C4067 XA4/XA4/A XA4/XA4/MN2/a_324_n18# 0.15fF
C4068 XA8/XA12/A VREF 0.02fF
C4069 XA2/DONE XA2/XA9/B 0.03fF
C4070 XA4/CN0 XA1/CN1 0.06fF
C4071 XA2/CP0 XA2/XA5/MN3/a_324_n18# 0.15fF
C4072 AVDD XA6/XA1/XA1/MP3/S 0.14fF
C4073 XA5/XA9/Y AVSS 0.22fF
C4074 D<4> XA4/CN1 0.42fF
C4075 XA5/XA5/MN1/a_324_n18# XA5/XA5/MN0/a_324_n18# 0.01fF
C4076 D<6> AVSS 2.30fF
C4077 XA1/XA1/XA5/MN2/S XA20/CNO 0.01fF
C4078 XA0/XA4/A AVSS 1.03fF
C4079 XA20/CPO XA2/XA1/XA1/MP3/G 0.14fF
C4080 XA0/CP0 XA3/CN1 0.14fF
C4081 XA5/XA4/A XA5/XA1/XA2/Y 0.19fF
C4082 XA2/XA11/MP0/a_216_n18# XA2/XA11/A 0.07fF
C4083 XA5/CN0 XA1/CN1 0.05fF
C4084 XA8/XA1/XA0/MN1/a_324_n18# XA8/XA1/XA1/MN0/a_324_n18# 0.01fF
C4085 XA2/XA1/XA1/MP2/a_216_n18# XA2/XA1/XA1/MP3/a_216_n18# 0.01fF
C4086 XA5/XA3/MN1/a_324_n18# XA5/CN1 0.16fF
C4087 XA0/XA6/MP3/a_216_n18# AVDD 0.08fF
C4088 XA8/XA8/MP0/a_216_n18# AVDD 0.09fF
C4089 VREF XA2/XA1/XA5/MP2/S 0.03fF
C4090 XA5/XA9/MN1/a_324_n18# XA5/XA9/A 0.07fF
C4091 XDAC2/XC1/XRES8/B XDAC2/XC1/XRES1A/B 0.12fF
C4092 XA8/EN XA7/XA6/MP3/S 0.02fF
C4093 XA0/XA2/MP3/a_216_n18# D<8> 0.02fF
C4094 XA8/EN XA7/XA7/MP0/a_216_n18# 0.07fF
C4095 XA6/XA3/MP2/a_216_n18# D<2> 0.01fF
C4096 D<1> XA7/XA1/XA2/Y 0.02fF
C4097 XA6/EN D<4> 0.02fF
C4098 XA3/XA1/XA1/MN2/a_324_n18# XA4/EN 0.01fF
C4099 XA4/XA1/XA2/Y XA20/CNO 0.22fF
C4100 XA2/EN XA2/XA2/MN0/a_324_n18# 0.07fF
C4101 XA4/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C4102 XA8/EN XA7/CN1 0.10fF
C4103 XA7/XA8/MP0/a_216_n18# XA7/XA9/MP0/a_216_n18# 0.01fF
C4104 XA5/XA11/A AVSS 0.27fF
C4105 XA5/CP0 XA5/EN 0.03fF
C4106 VREF XA1/EN 1.22fF
C4107 XA5/XA9/Y XA5/XA9/B 0.15fF
C4108 XA8/EN XA8/ENO 0.05fF
C4109 D<2> XA0/CP0 0.05fF
C4110 XA2/XA9/B D<6> 0.05fF
C4111 XA3/XA2/MP1/a_216_n18# VREF 0.02fF
C4112 XA20/XA2/MN6/a_324_n18# XA20/XA3/CO 0.08fF
C4113 XA7/XA3/MN2/a_324_n18# AVSS 0.01fF
C4114 XA4/XA6/MP3/S D<4> 0.02fF
C4115 XA20/XA4/MP0/S XA20/XA3/CO 0.10fF
C4116 XA0/XA9/Y XA0/CEO 0.01fF
C4117 XA5/XA1/XA5/MP1/S EN 0.03fF
C4118 D<2> XA6/XA6/MN1/S 0.01fF
C4119 XB2/XA3/B XB2/XA3/MP0/S 0.11fF
C4120 XA2/EN XA2/XA1/XA4/MN2/a_324_n18# 0.08fF
C4121 XA5/XA2/MN0/a_324_n18# AVSS 0.01fF
C4122 XA3/XA1/XA4/MN1/S AVDD 0.02fF
C4123 XA8/XA1/XA1/MP2/a_216_n18# XA8/XA1/XA1/MP3/G 0.01fF
C4124 XA4/XA2/A XA4/XA1/XA5/MP2/S 0.06fF
C4125 XA8/CN0 XA8/XA6/MP1/a_216_n18# 0.15fF
C4126 XA2/XA2/MP3/a_216_n18# AVDD 0.07fF
C4127 XA4/XA6/MN2/a_324_n18# XA4/XA6/MN3/a_324_n18# 0.01fF
C4128 XA5/CN1 EN 0.02fF
C4129 XDAC1/XC0/XRES4/B XDAC1/XC0/XRES16/B 0.25fF
C4130 XB2/XA3/MP0/S AVSS 0.22fF
C4131 XA3/XA5/MN3/a_324_n18# XA3/CN0 0.01fF
C4132 XA5/XA9/B XA5/XA11/A 0.02fF
C4133 XA1/XA6/MN1/a_324_n18# XA1/XA6/MN2/a_324_n18# 0.01fF
C4134 XA5/CN1 XA5/XA3/MN0/a_324_n18# 0.10fF
C4135 XA2/XA6/MN2/a_324_n18# XA2/XA6/MN3/a_324_n18# 0.01fF
C4136 SARP AVSS 111.47fF
C4137 XA1/EN XA0/XA7/MP0/a_216_n18# 0.07fF
C4138 XA7/XA12/A XA6/CEO 0.18fF
C4139 XA0/CP0 D<3> 0.05fF
C4140 XA20/XA2a/MN3/a_324_n18# XA20/XA3/CO 0.15fF
C4141 XA5/EN XA4/XA1/XA1/MN3/a_324_n18# 0.01fF
C4142 XA20/XA3/N2 XA20/XA3/CO 0.21fF
C4143 D<3> XA5/XA6/MP1/S 0.02fF
C4144 XDAC1/XC64b<1>/XRES1A/B XDAC1/X16ab/XRES4/B 0.01fF
C4145 XA3/XA3/MP0/a_216_n18# AVDD 0.08fF
C4146 XDAC1/XC32a<0>/XRES4/B XDAC1/XC128a<1>/XRES16/B 0.03fF
C4147 XB1/XA4/MN1/a_324_334# AVSS 0.01fF
C4148 XA0/XA1/XA0/MP1/a_216_n18# XA0/XA1/XA1/MP0/a_216_n18# 0.01fF
C4149 XA4/EN XA3/XA1/XA1/MP2/a_216_n18# 0.02fF
C4150 XA2/EN XA1/XA1/XA1/MN2/a_324_n18# 0.01fF
C4151 XA4/XA1/XA5/MP0/a_216_n18# EN 0.16fF
C4152 XDAC1/X16ab/XRES1B/B SARP 1.79fF
C4153 XA6/XA1/XA5/MN2/a_324_n18# XA6/XA1/XA5/MN1/a_324_n18# 0.01fF
C4154 XA20/CPO XA3/XA4/A 0.03fF
C4155 EN XA0/XA1/XA4/MP1/S 0.03fF
C4156 D<6> CK_SAMPLE 0.10fF
C4157 XA20/XA3/CO XA8/CP0 0.02fF
C4158 XB2/XA3/MP2/a_216_n18# XB2/XA4/GNG 0.02fF
C4159 XA8/XA2/MN2/a_324_n18# AVSS 0.01fF
C4160 XB1/M4/G XB1/XA3/MP0/S 0.03fF
C4161 XA0/XA6/MN3/S AVSS 0.13fF
C4162 XA1/XA1/XA2/Y XA1/CN0 0.02fF
C4163 XA6/CN0 XA20/CPO 0.06fF
C4164 XA5/XA3/MP0/a_216_n18# XA5/XA2/A 0.08fF
C4165 XA2/XA1/XA2/Y XA2/XA1/XA4/MN0/a_324_n18# 0.02fF
C4166 XDAC1/XC128a<1>/XRES16/B XDAC1/XC128a<1>/XRES4/B 0.25fF
C4167 XA4/XA4/A XA3/CN1 0.07fF
C4168 XA8/ENO D<0> 0.36fF
C4169 XA1/XA9/Y AVDD 0.58fF
C4170 XA3/XA1/XA5/MP2/S VREF 0.03fF
C4171 XA5/XA2/MP1/a_216_n18# VREF 0.02fF
C4172 XA3/XA13/MP1/a_216_334# AVDD 0.17fF
C4173 D<6> EN 0.05fF
C4174 XA5/XA2/MP2/a_216_n18# XA5/XA2/MP3/a_216_n18# 0.01fF
C4175 XA0/XA4/A EN 0.23fF
C4176 XA8/XA1/XA5/MN2/S AVDD 0.02fF
C4177 XDAC2/XC64a<0>/XRES16/B XDAC2/XC32a<0>/XRES16/B 0.41fF
C4178 XA7/XA3/MP2/a_216_n18# AVDD 0.07fF
C4179 XA0/CP1 D<4> 0.05fF
C4180 XA5/XA9/A AVDD 0.62fF
C4181 XA2/XA4/MN0/a_324_n18# AVSS 0.01fF
C4182 XA6/XA1/XA2/Y XA20/CPO 0.22fF
C4183 XA7/EN AVSS 1.21fF
C4184 XA0/XA6/MN2/a_324_n18# XA0/XA6/MN1/a_324_n18# 0.01fF
C4185 XA7/XA1/XA2/Y XA7/CN0 0.03fF
C4186 XA2/XA2/A VREF 0.36fF
C4187 XA20/XA3/N1 XA20/XA2/MN3/a_324_n18# 0.02fF
C4188 XDAC2/XC64b<1>/XRES16/B XDAC2/X16ab/XRES4/B 0.03fF
C4189 XA8/XA9/MP1/a_216_334# AVDD 0.09fF
C4190 XB2/XCAPB1/XCAPB0/m3_324_308# XB2/XA4/GNG 0.07fF
C4191 XA2/XA9/B XA2/XA6/MP1/S 0.07fF
C4192 XA5/EN XA20/CNO 0.93fF
C4193 XA5/CEO AVSS 0.69fF
C4194 AVDD XB1/XA3/MP0/S 0.23fF
C4195 XA1/CP0 XDAC1/X16ab/XRES16/B 0.01fF
C4196 XA1/XA4/MP2/a_216_n18# VREF 0.03fF
C4197 XA3/XA1/XA5/MP1/S VREF 0.02fF
C4198 XA8/XA1/XA4/MN1/S AVDD 0.02fF
C4199 XA7/XA1/XA1/MP1/a_216_n18# AVDD 0.07fF
C4200 XDAC2/XC128b<2>/XRES8/B XDAC2/XC128b<2>/XRES16/B 1.42fF
C4201 XA6/XA2/A D<2> 0.07fF
C4202 XA6/XA9/B XA6/XA6/MN3/S 0.09fF
C4203 XA6/XA9/A AVDD 0.62fF
C4204 XA2/XA5/MP0/a_216_n18# AVDD 0.08fF
C4205 XA7/XA1/XA1/MP0/a_216_n18# XA7/XA1/XA1/MP1/a_216_n18# 0.01fF
C4206 XA3/XA1/XA4/MP2/S EN 0.03fF
C4207 XA0/XA11/A AVSS 0.27fF
C4208 XA4/DONE XA4/XA9/A 0.07fF
C4209 XA1/XA1/XA1/MP0/a_216_n18# AVDD 0.14fF
C4210 XA2/XA1/XA4/MN1/S XA2/XA1/XA4/MN2/S 0.04fF
C4211 VREF XA0/XA2/MP2/a_216_n18# 0.03fF
C4212 XA1/XA9/Y XA1/XA9/MN1/S 0.12fF
C4213 D<3> XA4/XA4/A 0.01fF
C4214 XA5/XA4/A XA5/XA1/XA4/MN1/S 0.02fF
C4215 D<0> XA8/CN0 0.40fF
C4216 XA2/CP0 XA0/CP1 0.07fF
C4217 XA3/XA12/MP0/a_216_n18# XA3/XA12/A 0.07fF
C4218 AVDD XA2/XA1/XA2/Y 0.33fF
C4219 XA4/EN XA3/XA1/XA2/MP0/a_216_n18# 0.08fF
C4220 XA4/XA7/MN0/a_324_n18# XA4/XA9/B 0.01fF
C4221 XA5/XA9/B XA5/CEO 0.03fF
C4222 XA1/XA4/MN2/a_324_n18# XA1/XA4/MN1/a_324_n18# 0.01fF
C4223 D<6> XA2/XA7/MP0/a_216_n18# 0.08fF
C4224 XA8/EN XA7/XA1/XA1/MN3/a_324_n18# 0.02fF
C4225 XDAC1/XC0/XRES2/B SARP 3.05fF
C4226 XA4/CP0 XA4/XA4/MN1/a_324_n18# 0.03fF
C4227 XA2/XA12/MN0/a_324_n18# XA2/XA13/MN1/a_324_n18# 0.01fF
C4228 XA1/CN0 D<8> 0.13fF
C4229 XA0/XA6/MN3/S CK_SAMPLE 0.02fF
C4230 XA2/XA1/XA1/MP3/S XA2/XA1/XA1/MP3/G 0.04fF
C4231 XA20/XA2/MP0/a_216_n18# AVDD 0.17fF
C4232 XA8/XA3/MP1/a_216_n18# VREF 0.02fF
C4233 XA0/XA3/MN0/a_324_n18# D<8> 0.10fF
C4234 XA8/XA11/A XA8/CEO 0.01fF
C4235 XA6/XA1/XA5/MN2/a_324_n18# XA6/XA2/MN0/a_324_n18# 0.01fF
C4236 XA0/CEO XA0/CEIN 0.04fF
C4237 XA3/CN0 XA3/XA9/B 0.07fF
C4238 XA6/XA9/Y XA5/CEO 0.01fF
C4239 XA2/CP0 XA2/XA6/MP0/a_216_n18# 0.08fF
C4240 XA2/EN XA2/XA1/XA1/MN1/a_324_n18# 0.08fF
C4241 XA2/XA6/MP1/S CK_SAMPLE 0.03fF
C4242 XA3/XA2/MP1/a_216_n18# XA3/XA2/A 0.15fF
C4243 XA0/XA4/A XA0/XA4/MN2/a_324_n18# 0.15fF
C4244 XA5/XA4/MP1/a_216_n18# XA5/XA4/A 0.15fF
C4245 XB2/XA3/B XB2/XCAPB1/XCAPB4/m3_9756_132# 0.07fF
C4246 XA20/XA1/MN0/a_324_n18# XA20/XA9/A 0.08fF
C4247 XA3/XA2/MP3/a_216_n18# XA3/CN1 0.02fF
C4248 XA6/XA9/B XA6/XA9/MN1/S 0.02fF
C4249 XA20/XA1/MP0/S AVDD 0.58fF
C4250 XA1/XA2/MP2/a_216_n18# AVDD 0.07fF
C4251 XA1/XA2/A XA1/XA2/MN2/a_324_n18# 0.15fF
C4252 XA3/CP0 XA20/CPO 0.06fF
C4253 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC128a<1>/XRES1A/B 0.63fF
C4254 XDAC1/XC1/XRES16/B XDAC1/XC1/XRES1A/B 1.60fF
C4255 XA7/EN CK_SAMPLE 0.09fF
C4256 XA4/XA4/A XA4/XA4/MP3/a_216_n18# 0.15fF
C4257 XA20/CNO XA7/XA2/A 0.04fF
C4258 XA7/XA5/MP3/a_216_n18# AVDD 0.07fF
C4259 XDAC2/XC64a<0>/XRES4/B SARN 6.32fF
C4260 XA7/EN XA6/XA1/XA1/MP1/a_216_n18# 0.01fF
C4261 XA8/XA4/MP0/a_216_n18# VREF 0.02fF
C4262 XA1/CP0 XA1/XA5/MP0/a_216_n18# 0.07fF
C4263 XA5/XA3/MP0/a_216_n18# XA5/CN1 0.07fF
C4264 XA4/XA1/XA2/Y XA4/XA1/XA5/MN2/a_324_n18# 0.07fF
C4265 XA0/XA1/XA5/MP1/S XA0/XA1/XA5/MP2/S 0.04fF
C4266 XB2/M3/a_324_n18# XB2/M4/a_324_n18# 0.01fF
C4267 XDAC1/XC128b<2>/XRES4/B XDAC1/X16ab/XRES8/B 0.01fF
C4268 XA4/XA9/B XA4/XA8/MN0/a_324_n18# 0.01fF
C4269 XA7/XA9/MN1/S AVDD 0.01fF
C4270 XDAC1/XC128a<1>/XRES1A/B XDAC1/XC128a<1>/XRES1B/B 0.01fF
C4271 XA0/CP0 XDAC1/XC1/XRES16/B 0.20fF
C4272 XA2/XA13/MP1/a_216_n18# XA2/CEO 0.01fF
C4273 XA7/EN EN 1.03fF
C4274 XDAC2/X16ab/XRES16/B AVSS 16.03fF
C4275 XA8/EN XA7/XA1/XA2/Y 0.14fF
C4276 XA3/CN0 XA1/CN1 0.08fF
C4277 XA4/XA9/B AVSS 0.61fF
C4278 XA7/XA4/MN1/a_324_n18# XA7/XA4/MN0/a_324_n18# 0.01fF
C4279 XB1/XCAPB1/XCAPB0/m3_9756_132# XB1/XA3/B 0.07fF
C4280 XB1/XCAPB1/XCAPB4/m3_9828_132# XB1/XA4/GNG 0.03fF
C4281 XA2/XA3/MP1/a_216_n18# AVDD 0.07fF
C4282 XA1/XA9/MP1/a_216_n18# AVDD 0.09fF
C4283 XA3/XA11/MP0/a_216_n18# XA3/XA9/MP1/a_216_334# 0.01fF
C4284 XA6/XA9/B XA6/XA9/MP1/a_216_n18# 0.07fF
C4285 XA1/XA11/MP1/a_216_n18# XA0/CEO 0.07fF
C4286 XA7/XA11/MP1/S AVDD 0.18fF
C4287 XA5/XA3/MP1/a_216_n18# AVDD 0.07fF
C4288 XA0/XA5/MP2/a_216_n18# VREF 0.03fF
C4289 XDAC2/X16ab/XRES4/B SARN 6.32fF
C4290 XA4/CN0 AVSS 1.00fF
C4291 XA4/CEO XA4/XA12/A 0.10fF
C4292 XA4/XA1/XA4/MP2/S AVDD 0.11fF
C4293 XA8/XA5/MN2/a_324_n18# XA8/XA5/MN3/a_324_n18# 0.01fF
C4294 XA8/XA1/XA5/MP2/S XA8/XA4/A 0.02fF
C4295 XA2/CN1 XA0/CN0 0.16fF
C4296 XA6/XA1/XA1/MN1/a_324_n18# XA20/CNO 0.07fF
C4297 XA20/XA1/MN6/a_324_n18# SARP 0.08fF
C4298 XA3/XA2/A XA3/XA1/XA5/MP2/S 0.06fF
C4299 XA0/XA5/MN3/a_324_n18# XA0/XA5/MN2/a_324_n18# 0.01fF
C4300 XA6/XA2/A XA8/EN 0.03fF
C4301 XA2/XA4/A XA3/EN 0.11fF
C4302 XA1/XA9/Y XA1/XA9/A 0.04fF
C4303 XA1/XA2/A XA20/CNO 0.04fF
C4304 XA3/CN0 XA3/XA6/MP1/a_216_n18# 0.15fF
C4305 XB1/XA4/GNG XB1/XA1/Y 0.03fF
C4306 XA5/CN0 AVSS 1.14fF
C4307 XA0/XA9/A XA0/XA8/MP0/a_216_n18# 0.07fF
C4308 XA4/XA6/MN3/S XA4/XA9/B 0.09fF
C4309 XB1/CKN XB1/XA4/GNG 0.25fF
C4310 XA4/XA3/MP3/a_216_n18# XA4/CN1 0.15fF
C4311 XA8/XA2/MN1/a_324_n18# XA8/XA2/MN0/a_324_n18# 0.01fF
C4312 XA7/XA6/MP1/S VREF 0.04fF
C4313 XA1/CP0 XA1/XA4/MP3/a_216_n18# 0.02fF
C4314 XA8/XA2/MN2/a_324_n18# XA8/CN1 0.02fF
C4315 XA4/XA4/MN0/a_324_n18# AVSS 0.01fF
C4316 XA6/EN XA4/XA1/XA1/MP3/G 0.01fF
C4317 XA3/XA2/A XA2/XA2/A 0.03fF
C4318 XA4/XA3/MP0/a_216_n18# XA4/XA2/MP3/a_216_n18# 0.01fF
C4319 XA5/XA4/MP1/a_216_n18# VREF 0.02fF
C4320 XA0/XA1/XA4/MP0/a_216_n18# XA1/EN 0.08fF
C4321 XA6/XA5/MP1/a_216_n18# VREF 0.02fF
C4322 XB1/XA7/MP1/a_216_334# XB1/XA2/MP0/G 0.07fF
C4323 XA8/XA2/MP3/a_216_n18# XA8/CN1 0.02fF
C4324 XA4/XA1/XA5/MN1/S XA20/CNO 0.01fF
C4325 XA5/XA2/A XA5/XA4/A 0.14fF
C4326 XA7/XA9/MP0/a_216_n18# XA7/XA9/A 0.14fF
C4327 XA5/XA9/Y XA5/DONE 0.06fF
C4328 XA5/XA1/XA1/MP3/a_216_n18# XA5/XA1/XA1/MP2/a_216_n18# 0.01fF
C4329 XA6/XA7/MN0/a_324_n18# XA7/EN 0.08fF
C4330 XA2/XA9/MN0/a_324_n18# XA2/XA9/MN1/a_324_n18# 0.01fF
C4331 XA5/XA9/B XA5/CN0 0.07fF
C4332 D<2> XA6/XA6/MP1/S 0.02fF
C4333 XA4/XA1/XA1/MN1/a_324_n18# XA20/CNO 0.07fF
C4334 XA3/XA6/MP3/S XA4/EN 0.02fF
C4335 XA6/XA11/MP1/S VREF 0.01fF
C4336 XA20/XA12/Y DONE 0.07fF
C4337 XA0/XA9/MN1/S XA0/XA9/Y 0.12fF
C4338 DONE AVSS 0.31fF
C4339 XA1/XA1/XA5/MN0/a_324_n18# XA1/XA1/XA4/MN2/a_324_n18# 0.01fF
C4340 XA5/XA1/XA5/MP1/a_216_n18# XA5/XA1/XA5/MP2/a_216_n18# 0.01fF
C4341 XA2/XA3/MP3/a_216_n18# XA2/CN1 0.15fF
C4342 XA20/XA3/N1 XA20/XA2/MN5/a_324_n18# 0.02fF
C4343 XDAC1/X16ab/XRES1A/B SARP 1.50fF
C4344 XA2/EN XA0/XA2/A 0.03fF
C4345 XA8/ENO XA8/CN0 0.06fF
C4346 D<4> XA4/EN 0.03fF
C4347 XDAC2/XC64a<0>/XRES1A/B XDAC2/XC64a<0>/XRES2/B 0.25fF
C4348 XA1/EN XA0/XA1/XA1/MP3/S 0.10fF
C4349 XA3/CN0 XA3/XA1/XA1/MP3/G 0.02fF
C4350 XA4/XA3/MN2/a_324_n18# AVSS 0.01fF
C4351 XA2/XA3/MP0/a_216_n18# XA2/XA2/MP3/a_216_n18# 0.01fF
C4352 XA4/XA11/A XA4/CEO 0.01fF
C4353 XA7/XA5/MP0/a_216_n18# XA7/XA5/MP1/a_216_n18# 0.01fF
C4354 XB2/XA4/GNG XDAC2/XC1/XRES2/B 0.19fF
C4355 XA4/XA9/B CK_SAMPLE 0.09fF
C4356 XA7/XA5/MN2/a_324_n18# AVSS 0.01fF
C4357 XA6/CN1 XA6/XA3/MN3/a_324_n18# 0.15fF
C4358 XA4/XA6/MN1/S XA4/XA9/B 0.05fF
C4359 XB1/XCAPB1/XCAPB2/m3_324_308# XB1/XA4/GNG 0.07fF
C4360 XA0/XA3/MP3/a_216_n18# VREF 0.03fF
C4361 VREF XA0/XA3/MP2/a_216_n18# 0.03fF
C4362 XDAC1/XC32a<0>/XRES16/B XDAC1/XC64a<0>/XRES16/B 0.41fF
C4363 AVDD XB1/XA5/MP1/a_216_n18# 0.13fF
C4364 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128a<1>/XRES4/B 0.01fF
C4365 XA6/XA9/A XA6/XA9/MN0/a_324_n18# 0.15fF
C4366 XA8/XA12/A XA8/XA11/MN1/a_324_n18# 0.01fF
C4367 XA20/XA3/MP1/a_216_n18# XA20/XA3a/A 0.01fF
C4368 XB2/XA4/MN1/S AVDD 0.01fF
C4369 XA4/CN0 CK_SAMPLE 0.09fF
C4370 D<7> XA0/CN0 0.06fF
C4371 XDAC1/XC128b<2>/XRES8/B SARP 11.94fF
C4372 XB1/XCAPB1/XCAPB0/m3_252_308# XB1/XA3/B 0.02fF
C4373 SAR_IP SARP 1.07fF
C4374 XB2/XA3/B XDAC2/XC1/XRES8/B 0.06fF
C4375 XA2/CN0 D<4> 0.07fF
C4376 XA6/XA1/XA5/MN2/a_324_n18# XA6/XA1/XA2/Y 0.07fF
C4377 XA6/XA12/A XA6/XA11/A 0.07fF
C4378 XA4/CN1 XA4/XA3/MN3/a_324_n18# 0.15fF
C4379 XB1/M2/a_324_n18# XB1/M4/G 0.15fF
C4380 XA6/XA1/XA1/MP0/a_216_n18# AVDD 0.15fF
C4381 XA5/CN0 CK_SAMPLE 0.07fF
C4382 XA8/XA1/XA1/MN2/a_324_n18# XA8/XA1/XA1/MN3/a_324_n18# 0.01fF
C4383 XA2/CP0 XA4/EN 0.04fF
C4384 XA7/XA4/A VREF 0.37fF
C4385 AVDD XA8/XA5/MP1/a_216_n18# 0.07fF
C4386 XA1/CP0 XA1/XA6/MP0/a_216_n18# 0.08fF
C4387 XDAC2/XC1/XRES8/B AVSS 9.01fF
C4388 XA6/CEO XA6/XA12/A 0.11fF
C4389 XA4/XA3/MP2/a_216_n18# D<4> 0.01fF
C4390 XA4/CN0 EN 0.07fF
C4391 XA1/XA2/MN2/a_324_n18# XA1/CN1 0.02fF
C4392 XA8/XA2/MP1/a_216_n18# XA8/CN1 0.01fF
C4393 XA6/CP0 AVSS 0.91fF
C4394 XA3/XA1/XA5/MN1/a_324_n18# XA3/XA1/XA2/Y 0.08fF
C4395 XA5/XA1/XA1/MP3/a_216_n18# XA20/CPO 0.08fF
C4396 XA7/XA4/MN2/a_324_n18# XA7/CP0 0.01fF
C4397 XA20/CPO XA20/XA3/CO 0.29fF
C4398 XA1/XA12/A VREF 0.03fF
C4399 XA5/CEO XA6/XA12/MP0/a_216_n18# 0.08fF
C4400 XA0/XA8/MP0/a_216_n18# AVDD 0.09fF
C4401 XA20/CNO XA3/XA1/XA1/MN1/a_324_n18# 0.07fF
C4402 XA0/CP1 XA1/CN0 0.01fF
C4403 XA20/XA3/MP0/a_216_n18# XA20/XA3a/MP3/a_216_n18# 0.01fF
C4404 XA1/CP0 XA3/CP0 0.16fF
C4405 XA5/CN0 EN 0.06fF
C4406 XA8/XA4/A AVDD 1.49fF
C4407 XA5/XA2/A VREF 0.36fF
C4408 XA6/XA3/MP0/a_216_n18# XA6/XA2/A 0.08fF
C4409 XA6/XA2/MP1/a_216_n18# XA6/XA2/MP2/a_216_n18# 0.01fF
C4410 XA5/XA1/XA5/MN2/S AVDD 0.02fF
C4411 D<4> SARN 0.03fF
C4412 XA5/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C4413 XA6/XA1/XA4/MN2/S XA6/XA1/XA4/MN1/S 0.04fF
C4414 XA3/XA4/MN2/a_324_n18# AVSS 0.01fF
C4415 XA3/XA11/MP1/S VREF 0.01fF
C4416 XA1/XA1/XA4/MN1/S XA1/EN 0.02fF
C4417 D<6> XA2/CN1 0.83fF
C4418 XA2/CP0 XA2/CN0 3.92fF
C4419 XA6/XA2/MP1/a_216_n18# AVDD 0.08fF
C4420 DONE CK_SAMPLE 0.26fF
C4421 XA6/XA3/MP3/a_216_n18# D<2> 0.02fF
C4422 XA20/XA3/N1 XA20/XA3/CO 0.30fF
C4423 XA5/EN XA4/XA1/XA4/MP2/S 0.02fF
C4424 XA5/XA4/A XA5/XA1/XA5/MP1/S 0.02fF
C4425 XA3/XA2/MN2/a_324_n18# XA3/XA2/MN3/a_324_n18# 0.01fF
C4426 XA1/XA9/MP1/a_216_n18# XA1/XA9/A 0.08fF
C4427 XA6/XA12/MN0/a_324_n18# XA6/XA11/MN1/a_324_n18# 0.01fF
C4428 XA1/XA1/XA1/MN0/a_324_n18# XA1/XA1/XA0/MN1/a_324_n18# 0.01fF
C4429 XA20/XA12/Y XA20/XA10/MN1/a_324_n18# 0.08fF
C4430 XA4/XA6/MP3/a_216_n18# D<4> 0.15fF
C4431 XA1/CEO XA1/XA9/B 0.03fF
C4432 XA5/XA13/MP1/a_216_334# AVDD 0.17fF
C4433 XA2/XA1/XA0/MN1/a_324_n18# XA2/XA1/XA1/MN0/a_324_n18# 0.01fF
C4434 XA2/EN XA1/XA1/XA1/MN2/S 0.12fF
C4435 XA20/XA2a/MN2/a_324_n18# XA20/XA3/CO 0.15fF
C4436 XA1/XA11/A AVSS 0.27fF
C4437 XA8/XA1/XA1/MP2/S XA8/XA1/XA1/MP3/S 0.04fF
C4438 XA6/XA6/MP0/a_216_n18# XA6/XA5/MP3/a_216_n18# 0.01fF
C4439 XA5/CN1 XA5/XA4/A 0.58fF
C4440 XA2/XA9/A AVDD 0.62fF
C4441 XA1/CN0 XA1/XA5/MN3/a_324_n18# 0.01fF
C4442 XA20/XA4/MN5/a_324_n18# XA20/XA4/MN4/a_324_n18# 0.01fF
C4443 XDAC2/XC128a<1>/XRES8/B AVSS 9.08fF
C4444 XA6/XA6/MP3/S VREF 0.02fF
C4445 XA4/XA9/B XA4/XA9/A 0.29fF
C4446 XDAC1/X16ab/XRES8/B AVSS 9.08fF
C4447 XA2/CP0 SARN 0.03fF
C4448 XA7/XA9/B XA7/XA7/MN0/a_324_n18# 0.01fF
C4449 XA20/CNO XA1/CN1 0.20fF
C4450 XB2/XA4/GNG XB2/XCAPB1/XCAPB3/m3_9828_132# 0.04fF
C4451 VREF XA0/CN0 0.69fF
C4452 XDAC1/XC64a<0>/XRES8/B XDAC1/XC64a<0>/XRES1B/B 0.12fF
C4453 XA7/XA2/MN0/a_324_n18# AVSS 0.01fF
C4454 XA20/XA3/MN2/a_324_n18# SARN 0.15fF
C4455 XA20/XA3a/MN2/a_324_n18# XA20/XA3a/A 0.15fF
C4456 XA3/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C4457 XDAC2/XC32a<0>/XRES2/B XDAC2/XC32a<0>/XRES1B/B 0.23fF
C4458 XDAC1/XC32a<0>/C1A AVSS 0.01fF
C4459 XA8/XA3/MP3/a_216_n18# XA8/CN1 0.15fF
C4460 XA3/XA2/A XA3/XA1/XA2/Y 0.01fF
C4461 XA20/XA3/MN4/a_324_n18# XA20/XA3/MN3/a_324_n18# 0.01fF
C4462 XDAC2/XC128a<1>/XRES1B/B XDAC2/XC128a<1>/XRES8/B 0.12fF
C4463 XA3/XA11/A AVDD 0.45fF
C4464 AVSS XA8/XA6/MN1/S 0.16fF
C4465 XDAC2/XC128a<1>/XRES16/B XDAC2/XC32a<0>/XRES4/B 0.03fF
C4466 EN XA0/XA1/XA4/MP2/a_216_n18# 0.16fF
C4467 XDAC1/X16ab/XRES1B/B XDAC1/X16ab/XRES8/B 0.12fF
C4468 XA5/XA9/MN1/S AVSS 0.15fF
C4469 XA1/XA2/MP0/a_216_n18# EN 0.08fF
C4470 XA6/XA9/Y XA6/XA11/MP0/a_216_n18# 0.08fF
C4471 XA6/CP0 CK_SAMPLE 0.09fF
C4472 XA2/CN1 SARP 0.07fF
C4473 XB2/M4/G XB2/XA3/MP0/S 0.03fF
C4474 XDAC1/XC64b<1>/XRES16/B XDAC1/X16ab/XRES2/B 0.01fF
C4475 XA7/EN XA6/XA1/XA1/MP3/G 0.27fF
C4476 XA20/XA2/MN0/a_324_n18# SARP 0.02fF
C4477 XA8/XA9/MP0/a_216_n18# XA8/XA9/A 0.14fF
C4478 XA2/CP0 XA2/XA5/MP3/a_216_n18# 0.15fF
C4479 XA3/XA9/MP1/a_216_334# XA3/XA9/MP1/a_216_n18# 0.01fF
C4480 XDAC1/XC64b<1>/XRES8/B XDAC1/XC64b<1>/XRES16/B 1.42fF
C4481 XB2/M4/G SARP 0.05fF
C4482 XA3/XA11/A XA3/XA9/Y 0.14fF
C4483 XB1/XA1/MP0/G XB1/XA7/MN1/a_324_n18# 0.07fF
C4484 XA8/XA5/MN0/a_324_n18# XA8/XA4/A 0.07fF
C4485 XB1/XA4/MP1/a_216_n18# XB1/XA4/MP0/a_216_n18# 0.01fF
C4486 XA5/XA9/B XA5/XA9/MN1/S 0.02fF
C4487 XA0/XA4/MP1/a_216_n18# AVDD 0.07fF
C4488 XA7/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C4489 XA20/CPO XA1/EN 0.64fF
C4490 XA2/XA13/MP1/a_216_334# XA2/XA13/MP1/a_216_n18# 0.01fF
C4491 D<7> D<6> 1.47fF
C4492 XA1/XA2/MP2/a_216_n18# XA1/XA2/A 0.15fF
C4493 D<7> XA0/XA4/A 0.01fF
C4494 XDAC2/XC0/XRES16/B D<8> 0.22fF
C4495 XA5/XA1/XA5/MP2/S AVDD 0.08fF
C4496 XA7/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C4497 XA2/XA3/MP3/a_216_n18# VREF 0.03fF
C4498 XB1/M7/a_324_n18# SAR_IP 0.01fF
C4499 XA0/XA9/Y XA0/DONE 0.06fF
C4500 XA0/XA9/B AVSS 0.60fF
C4501 XDAC1/XC1/XRES4/B XDAC1/XC64a<0>/XRES8/B 0.01fF
C4502 XA5/XA1/XA5/MP1/S VREF 0.02fF
C4503 XA5/XA6/MP3/S AVDD 0.16fF
C4504 XA0/CEIN XB1/M8/a_324_334# 0.09fF
C4505 XA3/CN0 AVSS 0.89fF
C4506 XDAC1/XC32a<0>/XRES8/B XDAC1/XC32a<0>/XRES16/B 1.42fF
C4507 XA0/CEIN XB1/XA2/MP0/G 0.04fF
C4508 XA0/XA5/MP3/a_216_n18# VREF 0.02fF
C4509 XA2/XA4/A XA2/XA1/XA4/MP2/S 0.05fF
C4510 XA3/XA5/MP3/a_216_n18# VREF 0.02fF
C4511 XA2/XA6/MN1/S AVDD 0.01fF
C4512 XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MP3/a_216_n18# 0.07fF
C4513 XA2/XA3/MP1/a_216_n18# XA2/XA3/MP0/a_216_n18# 0.01fF
C4514 XA1/CEO XA2/XA12/MN0/a_324_n18# 0.07fF
C4515 XA5/CN1 VREF 0.76fF
C4516 XA20/CNO XA3/XA1/XA1/MP3/G 0.06fF
C4517 XA6/DONE AVDD 0.21fF
C4518 XA2/CN1 XA2/XA4/MN0/a_324_n18# 0.07fF
C4519 XA8/XA1/XA4/MN1/a_324_n18# XA8/XA1/XA4/MN2/a_324_n18# 0.01fF
C4520 XB1/XCAPB1/XCAPB4/m3_324_308# XB1/XA4/GNG 0.07fF
C4521 XDAC1/XC0/XRES4/B AVSS 5.40fF
C4522 XA8/XA1/XA2/Y XA8/XA1/XA5/MN1/a_324_n18# 0.09fF
C4523 XDAC2/XC64b<1>/XRES16/B XA1/CN0 0.01fF
C4524 XA2/XA1/XA4/MN0/a_324_n18# XA2/XA1/XA4/MN1/a_324_n18# 0.01fF
C4525 VREF XA1/XA5/MP1/a_216_n18# 0.02fF
C4526 XA7/XA8/MN0/a_324_n18# XA7/XA9/A 0.09fF
C4527 XA2/XA2/MN2/a_324_n18# XA2/XA2/MN3/a_324_n18# 0.01fF
C4528 CK_SAMPLE XA8/XA6/MN1/S 0.04fF
C4529 XA20/XA1/MN2/a_324_n18# XA20/XA1/MN3/a_324_n18# 0.01fF
C4530 XA6/XA12/MP0/a_216_n18# XA6/XA13/MP1/a_216_n18# 0.01fF
C4531 AVDD XA20/XA2a/MP1/a_216_n18# 0.09fF
C4532 XA0/XA1/XA5/MP1/S XA1/EN 0.02fF
C4533 AVDD XB1/XA0/MP0/a_216_n18# 0.15fF
C4534 XA8/CEO XA20/XA12/MP0/a_216_n18# 0.07fF
C4535 XA6/XA1/XA5/MP1/S XA6/XA4/A 0.02fF
C4536 XA6/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C4537 XA7/XA1/XA0/MN1/a_324_n18# XA7/XA1/XA1/MN0/a_324_n18# 0.01fF
C4538 XA0/XA4/MN0/a_324_n18# D<8> 0.07fF
C4539 D<7> SARP 0.28fF
C4540 XA0/XA3/MN2/a_324_n18# AVSS 0.01fF
C4541 XB1/XA4/GNG AVSS 5.21fF
C4542 XDAC1/XC64b<1>/XRES8/B XDAC1/XC0/XRES8/B 0.21fF
C4543 XB1/XCAPB1/XCAPB2/m3_9756_132# XB1/XA3/B 0.07fF
C4544 VREF XA3/XA4/MP3/a_216_n18# 0.03fF
C4545 XDAC1/XC32a<0>/XRES8/B XDAC1/XC32a<0>/XRES2/B 1.58fF
C4546 XA7/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C4547 XDAC1/XC64b<1>/XRES16/B XDAC1/XC0/XRES1A/B 0.04fF
C4548 XA5/XA1/XA2/Y XA20/CPO 0.23fF
C4549 XA7/XA7/MN0/a_324_n18# AVSS 0.01fF
C4550 XA20/XA2a/MP3/a_216_n18# XA20/XA2a/MP2/a_216_n18# 0.01fF
C4551 XA8/XA12/A XA8/XA11/MP1/S 0.06fF
C4552 XA6/XA1/XA4/MN1/S XA20/CPO 0.03fF
C4553 XA0/CEO XA0/XA12/A 0.11fF
C4554 XA2/CP0 XA2/XA5/MN2/a_324_n18# 0.15fF
C4555 XA20/XA2/MN1/a_324_n18# XA20/XA2/MN0/a_324_n18# 0.01fF
C4556 XB1/XA3/MP0/S XB1/XA1/Y 0.02fF
C4557 XA5/XA11/MP1/S AVDD 0.18fF
C4558 XA2/XA1/XA1/MP0/a_216_n18# XA2/XA1/XA1/MP1/a_216_n18# 0.01fF
C4559 XA5/XA9/Y VREF 0.03fF
C4560 XA6/XA9/MP0/a_216_n18# AVDD 0.09fF
C4561 D<6> VREF 1.73fF
C4562 XA6/XA1/XA1/MN3/a_324_n18# XA6/XA1/XA1/MP3/G 0.08fF
C4563 XA8/XA2/MP1/a_216_n18# XA8/XA2/MP0/a_216_n18# 0.01fF
C4564 XDAC2/XC64a<0>/XRES16/B AVSS 16.06fF
C4565 XA0/XA4/A VREF 0.37fF
C4566 XB1/CKN XB1/XA3/MP0/S 0.54fF
C4567 XA8/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C4568 XA8/CN0 XA8/XA5/MN3/a_324_n18# 0.01fF
C4569 XA7/XA1/XA5/MN1/a_324_n18# XA20/CNO 0.07fF
C4570 XA1/CP0 XDAC1/XC64a<0>/XRES16/B 0.16fF
C4571 XA5/CP0 AVSS 0.91fF
C4572 XA1/XA9/A XA2/XA9/A 0.02fF
C4573 XA0/XA9/B CK_SAMPLE 0.09fF
C4574 AVDD XB1/XA4/MP0/a_216_n18# 0.09fF
C4575 XA4/XA1/XA1/MP3/G XA4/EN 0.03fF
C4576 XA6/XA5/MP3/a_216_n18# AVDD 0.07fF
C4577 XA1/XA4/A XA1/XA1/XA5/MN1/S 0.02fF
C4578 XA3/CN0 CK_SAMPLE 0.09fF
C4579 XA1/CN0 XA1/XA5/MN1/a_324_n18# 0.02fF
C4580 XA5/XA11/A VREF 0.02fF
C4581 XA2/EN XA2/XA1/XA1/MP3/G 0.03fF
C4582 XA6/CN1 XA6/XA4/A 0.58fF
C4583 XA0/XA1/XA2/MN0/a_324_n18# XA0/XA1/XA1/MP3/G 0.06fF
C4584 XA5/XA9/MP1/a_216_n18# XA5/XA9/A 0.08fF
C4585 XA20/XA3a/MP0/a_216_n18# XA20/XA3/CO 0.08fF
C4586 D<7> XA1/XA4/MP0/a_216_n18# 0.01fF
C4587 XA3/XA11/MN1/a_324_n18# XA2/CEO 0.08fF
C4588 D<5> XA3/XA6/MP3/S 0.02fF
C4589 XA3/XA5/MN1/a_324_n18# XA3/CP0 0.15fF
C4590 XA3/XA5/MP1/a_216_n18# XA3/CP0 0.15fF
C4591 XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MP2/S 0.04fF
C4592 XA2/XA9/MN1/S AVDD 0.01fF
C4593 XA1/CN1 XA2/XA1/XA2/Y 0.02fF
C4594 XA8/XA11/MN1/a_324_n18# XA8/XA12/MN0/a_324_n18# 0.01fF
C4595 XA5/CEO XA6/XA11/MN1/a_324_n18# 0.08fF
C4596 XA20/XA9/MN0/a_324_334# XA20/XA11/Y 0.08fF
C4597 XA1/EN XA0/XA1/XA1/MP2/a_216_n18# 0.02fF
C4598 XA7/XA1/XA5/MN1/S AVSS 0.12fF
C4599 XA8/XA4/A XA7/XA2/A 0.03fF
C4600 XA2/CN0 XA1/CN0 0.57fF
C4601 XA3/XA1/XA4/MP0/a_216_n18# EN 0.07fF
C4602 XA3/CN0 EN 0.05fF
C4603 XA7/XA1/XA5/MP1/S EN 0.03fF
C4604 D<5> D<4> 0.28fF
C4605 XA1/XA1/XA2/Y XA1/XA1/XA4/MN2/S 0.05fF
C4606 XA7/XA1/XA5/MN2/S XA7/XA4/A 0.02fF
C4607 XDAC1/XC1/XRES8/B XDAC1/XC64a<0>/XRES1A/B 0.03fF
C4608 XA6/XA8/MN0/a_324_n18# XA7/EN 0.06fF
C4609 XA5/XA1/XA4/MN2/S AVDD 0.02fF
C4610 XA2/CN0 XA4/XA1/XA1/MP3/G 0.01fF
C4611 XA0/CP1 XA0/XA6/MP1/S 0.02fF
C4612 D<1> D<8> 0.18fF
C4613 XA1/XA12/A XA1/XA12/MN0/a_324_n18# 0.09fF
C4614 XA5/XA2/A XA4/XA2/A 0.03fF
C4615 XB1/M4/G XB1/M1/a_324_n18# 0.08fF
C4616 XA6/XA11/A AVDD 0.45fF
C4617 AVDD XA2/XA1/XA4/MN2/S 0.02fF
C4618 XA4/XA1/XA1/MN0/a_324_n18# XA4/XA1/XA0/MN1/a_324_n18# 0.01fF
C4619 EN XA5/XA1/XA5/MP0/a_216_n18# 0.16fF
C4620 XA3/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C4621 XA6/CN0 XA6/XA9/B 0.07fF
C4622 XA3/XA9/MN1/a_324_334# XA3/XA9/MN1/a_324_n18# 0.01fF
C4623 XA8/EN XA8/XA2/MN0/a_324_n18# 0.07fF
C4624 XA7/XA1/XA4/MN1/S XA7/XA4/A 0.02fF
C4625 XA6/CEO AVDD 1.64fF
C4626 XDAC1/XC0/XRES1A/B XDAC1/XC0/XRES8/B 0.12fF
C4627 XDAC1/XC0/XRES2/B XDAC1/XC0/XRES4/B 0.55fF
C4628 XA1/XA1/XA1/MP2/S AVDD 0.09fF
C4629 XA7/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C4630 XA4/EN XA3/EN 1.81fF
C4631 XA4/XA3/MP2/a_216_n18# XA4/XA3/MP3/a_216_n18# 0.01fF
C4632 XA6/XA9/MN1/a_324_n18# XA6/XA9/MN1/a_324_334# 0.01fF
C4633 XA4/CN0 XA2/CN1 0.31fF
C4634 SARN XA1/CN0 0.36fF
C4635 XA1/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C4636 XA4/XA12/MN0/a_324_n18# XA4/XA12/A 0.09fF
C4637 XA6/EN XA5/XA8/MP0/a_216_n18# 0.08fF
C4638 XA1/XA3/MN2/a_324_n18# XA1/CN1 0.16fF
C4639 XA3/CEO AVDD 0.74fF
C4640 XDAC1/XC32a<0>/XRES16/B XDAC1/XC64a<0>/XRES2/B 0.01fF
C4641 XA2/CP0 D<5> 3.01fF
C4642 XA8/EN XA8/XA1/XA4/MN2/a_324_n18# 0.08fF
C4643 XA1/CP0 XA1/EN 0.10fF
C4644 XA1/XA9/Y XA1/DONE 0.06fF
C4645 AVDD XA6/XA1/XA1/MN2/S 0.05fF
C4646 XA8/EN XA7/XA1/XA4/MN2/S 0.01fF
C4647 XA4/CP0 D<4> 0.23fF
C4648 XA5/CN0 XA2/CN1 0.07fF
C4649 XA8/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C4650 VREF XA1/XA5/MP3/a_216_n18# 0.02fF
C4651 XA1/XA5/MN0/a_324_n18# XA1/XA4/MN3/a_324_n18# 0.01fF
C4652 D<1> XA7/CP0 0.23fF
C4653 XA8/XA2/MP3/a_216_n18# VREF 0.02fF
C4654 XA5/CP0 CK_SAMPLE 0.08fF
C4655 XA2/XA6/MP1/S VREF 0.04fF
C4656 XA4/XA11/A XA4/XA12/A 0.07fF
C4657 XA3/CEO XA3/XA9/Y 0.03fF
C4658 XB2/XCAPB1/XCAPB0/m3_9828_132# XB2/XA4/GNG 0.03fF
C4659 XA1/XA5/MN2/a_324_n18# XA1/XA5/MN3/a_324_n18# 0.01fF
C4660 XA2/CN0 XA3/EN 0.33fF
C4661 XA3/XA1/XA4/MN0/a_324_n18# XA4/EN 0.07fF
C4662 XA5/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C4663 XDAC1/X16ab/XRES1A/B XDAC1/X16ab/XRES8/B 0.12fF
C4664 XA20/CPO XA2/XA1/XA2/MN0/a_324_n18# 0.01fF
C4665 XDAC1/XC128b<2>/XRES16/B XDAC1/XC128b<2>/XRES2/B 1.61fF
C4666 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128a<1>/XRES1A/B 0.12fF
C4667 XA4/XA3/MP1/a_216_n18# VREF 0.02fF
C4668 XA1/XA4/A XA1/XA3/MN3/a_324_n18# 0.01fF
C4669 XA1/XA4/MP0/a_216_n18# VREF 0.02fF
C4670 XA20/CNO AVSS 6.93fF
C4671 XA7/EN VREF 1.22fF
C4672 XA7/XA11/A XA6/CEO 0.09fF
C4673 XA20/XA0/MP1/a_216_n18# XA20/XA1/MP0/a_216_n18# 0.01fF
C4674 XA3/CN1 D<8> 2.16fF
C4675 XA6/XA1/XA1/MP3/S AVSS 0.02fF
C4676 XA4/XA1/XA5/MN1/a_324_n18# XA20/CNO 0.07fF
C4677 XA8/XA9/MP1/a_216_334# XA8/XA9/MP1/a_216_n18# 0.01fF
C4678 XDAC2/XC128b<2>/XRES8/B XDAC2/X16ab/XRES16/B 0.03fF
C4679 XDAC1/XC32a<0>/XRES2/B XDAC1/XC64a<0>/XRES2/B 0.05fF
C4680 XA5/CEO VREF 0.05fF
C4681 XA8/XA1/XA5/MN1/a_324_n18# XA8/XA1/XA5/MN2/a_324_n18# 0.01fF
C4682 XA5/XA1/XA1/MP3/G XA5/CN0 0.02fF
C4683 XA5/XA1/XA4/MN1/S XA20/CPO 0.04fF
C4684 XA8/XA1/XA4/MN1/a_324_n18# XA8/XA1/XA4/MN0/a_324_n18# 0.01fF
C4685 XDAC2/XC32a<0>/XRES1B/B XDAC2/XC32a<0>/XRES16/B 0.12fF
C4686 XA5/XA1/XA4/MP2/S AVDD 0.11fF
C4687 XDAC1/XC128b<2>/XRES8/B XDAC1/X16ab/XRES8/B 0.21fF
C4688 XA0/XA8/MP0/a_216_n18# XA0/XA9/MP0/a_216_n18# 0.01fF
C4689 XA5/XA1/XA1/MP3/G XA5/XA1/XA1/MP1/a_216_n18# 0.01fF
C4690 XA20/XA3/MP6/a_216_n18# AVDD 0.09fF
C4691 XA3/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C4692 XA2/XA3/MP2/a_216_n18# AVDD 0.07fF
C4693 VREF XA0/XA11/A 0.02fF
C4694 XDAC2/XC1/XRES4/B XDAC2/XC1/XRES2/B 0.55fF
C4695 XA7/XA1/XA5/MN1/S EN 0.01fF
C4696 D<2> D<8> 0.05fF
C4697 XA1/XA1/XA5/MP1/a_216_n18# XA1/XA1/XA5/MP0/a_216_n18# 0.01fF
C4698 XA1/XA1/XA1/MP1/a_216_n18# AVDD 0.07fF
C4699 XA7/XA1/XA1/MP2/S XA7/EN 0.01fF
C4700 XA7/CN0 D<8> 0.19fF
C4701 XB2/XCAPB1/XCAPB4/m3_252_308# XB2/XA3/B 0.02fF
C4702 XA20/XA2/MP4/a_216_n18# XA20/XA3/CO 0.07fF
C4703 XDAC1/XC64a<0>/XRES4/B AVSS 5.50fF
C4704 XA4/XA5/MP3/a_216_n18# VREF 0.02fF
C4705 XA8/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C4706 XA0/XA1/XA5/MP1/a_216_n18# XA0/XA1/XA5/MP0/a_216_n18# 0.01fF
C4707 XA20/CPO XA3/XA1/XA2/Y 0.24fF
C4708 XA7/XA1/XA4/MP2/S EN 0.03fF
C4709 XB2/CKN XB2/XA3/MN2/a_324_n18# 0.07fF
C4710 D<5> XA3/XA6/MP1/S 0.02fF
C4711 XA8/XA2/MP1/a_216_n18# VREF 0.02fF
C4712 XA1/XA9/B AVDD 0.79fF
C4713 XA3/XA4/MN3/a_324_n18# XA3/XA4/A 0.15fF
C4714 XA4/XA1/XA1/MP0/a_216_n18# XA4/XA1/XA0/MP1/a_216_n18# 0.01fF
C4715 XA8/XA1/XA1/MP3/G AVDD 0.65fF
C4716 XA20/XA2/MN6/a_324_n18# SARP 0.07fF
C4717 XA0/XA2/A XA0/XA1/XA5/MP2/S 0.06fF
C4718 XA5/CN0 XA5/XA4/A 0.12fF
C4719 XA7/XA3/MP1/a_216_n18# VREF 0.02fF
C4720 XA4/XA6/MP2/a_216_n18# XA4/CN0 0.08fF
C4721 XA6/XA1/XA5/MN2/S XA6/XA1/XA5/MN1/S 0.04fF
C4722 XB2/XA4/GNG XB2/XA4/MP1/a_216_n18# 0.02fF
C4723 D<3> D<8> 1.03fF
C4724 XA1/XA6/MP1/S CK_SAMPLE 0.03fF
C4725 XA8/XA1/XA5/MP2/S XA8/XA2/A 0.06fF
C4726 XA7/XA11/MP1/S XA7/CEO 0.02fF
C4727 XA1/XA6/MP2/a_216_n18# AVDD 0.09fF
C4728 XA3/XA1/XA4/MN1/S AVSS 0.10fF
C4729 XA3/XA1/XA5/MP2/a_216_n18# EN 0.16fF
C4730 AVDD XA2/XA11/MP1/S 0.19fF
C4731 XA8/XA1/XA2/Y XA7/EN 0.02fF
C4732 XA3/CEO XA4/XA12/MP0/a_216_n18# 0.08fF
C4733 XA8/XA1/XA4/MP2/a_216_n18# XA8/XA1/XA5/MP0/a_216_n18# 0.01fF
C4734 XA7/XA1/XA5/MP2/S AVDD 0.08fF
C4735 XB2/CKN XB2/XA3/MN0/a_324_n18# 0.09fF
C4736 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC64b<1>/XRES16/B 0.12fF
C4737 XA0/CP0 XA0/XA5/MP0/a_216_n18# 0.07fF
C4738 XA5/EN XA5/XA1/XA4/MN2/S 0.02fF
C4739 D<2> XA7/CP0 0.01fF
C4740 XA8/ENO XA8/XA7/MN0/a_324_n18# 0.08fF
C4741 XA0/XA4/MP0/a_216_n18# XA0/XA3/MP3/a_216_n18# 0.01fF
C4742 XA20/XA11/MN0/a_324_n18# XA20/XA12/Y 0.07fF
C4743 XDAC1/XC128b<2>/XRES1A/B SARP 1.50fF
C4744 XA0/XA1/XA4/MP2/S XA1/EN 0.02fF
C4745 XA4/CN1 XA3/CN1 0.12fF
C4746 XA20/CNO XA0/XA1/XA1/MN2/a_324_n18# 0.07fF
C4747 XA7/CN0 XA7/CP0 0.60fF
C4748 XA3/XA1/XA5/MN1/a_324_n18# XA3/XA1/XA5/MN0/a_324_n18# 0.01fF
C4749 XA8/XA4/MP2/a_216_n18# XA8/XA4/A 0.15fF
C4750 XA8/XA4/MN0/a_324_n18# AVSS 0.01fF
C4751 XA5/XA5/MP2/a_216_n18# XA5/CN0 0.01fF
C4752 XA2/XA1/XA1/MP3/G XA2/XA1/XA1/MN3/a_324_n18# 0.08fF
C4753 XDAC2/XC128b<2>/XRES1A/B XDAC2/X16ab/XRES1A/B 0.03fF
C4754 XA1/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C4755 XA6/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C4756 XA2/XA1/XA1/MP3/G XA2/XA1/XA2/MP0/a_216_n18# 0.08fF
C4757 XA7/XA4/MN0/a_324_n18# XA7/XA3/MN3/a_324_n18# 0.01fF
C4758 DONE XA8/XA9/B 0.05fF
C4759 XA7/XA1/XA5/MN0/a_324_n18# XA7/EN 0.07fF
C4760 XB2/XCAPB1/XCAPB2/m3_9756_132# XB2/XA3/B 0.07fF
C4761 XA1/XA9/B XA1/XA9/MN1/S 0.02fF
C4762 XA8/XA12/A XA8/XA9/Y 0.02fF
C4763 EN XA20/CNO 2.90fF
C4764 XA4/XA1/XA2/Y XA4/XA1/XA4/MN1/a_324_n18# 0.09fF
C4765 XA3/XA13/MP1/a_216_n18# AVDD 0.13fF
C4766 XA4/XA9/B VREF 0.12fF
C4767 AVDD XA8/XA6/MP2/a_216_n18# 0.09fF
C4768 XA1/XA9/Y AVSS 0.22fF
C4769 XA1/XA9/MN1/a_324_334# XA1/XA9/Y 0.09fF
C4770 XA7/XA4/MN0/a_324_n18# XA7/XA4/A 0.09fF
C4771 XA7/XA9/B XA7/XA9/MN1/S 0.02fF
C4772 XA8/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C4773 D<2> XA6/EN 0.03fF
C4774 XA20/CPO XA5/XA1/XA4/MP1/S 0.03fF
C4775 XA2/XA1/XA5/MP1/S XA2/XA1/XA5/MP2/S 0.04fF
C4776 XA7/XA4/A XA20/CPO 0.03fF
C4777 XA6/XA1/XA1/MP2/S XA7/EN 0.14fF
C4778 D<1> XA0/CP1 0.14fF
C4779 XA8/XA3/MP3/a_216_n18# VREF 0.02fF
C4780 XDAC2/XC0/XRES4/B AVSS 5.40fF
C4781 XA8/XA1/XA5/MN2/S AVSS 0.08fF
C4782 XA1/XA6/MN1/S AVDD 0.01fF
C4783 XA4/CN0 VREF 0.69fF
C4784 XA8/XA1/XA1/MN2/S XA20/CNO 0.03fF
C4785 XA6/XA1/XA2/Y XA6/XA1/XA5/MN1/a_324_n18# 0.09fF
C4786 XA5/XA9/A AVSS 0.31fF
C4787 XA2/XA6/MP0/a_216_n18# XA2/XA6/MP1/a_216_n18# 0.01fF
C4788 XA2/XA8/MN0/a_324_n18# XA2/XA9/A 0.09fF
C4789 XA7/CN0 XA6/EN 0.02fF
C4790 XDAC2/XC64b<1>/XRES16/B XDAC2/XC0/XRES16/B 0.41fF
C4791 XA1/XA1/XA4/MP1/S AVDD 0.14fF
C4792 D<3> XA4/CN1 0.01fF
C4793 XA8/XA4/MP1/a_216_n18# VREF 0.02fF
C4794 SAR_IP XB1/XA4/GNG 0.02fF
C4795 XA3/XA11/A XA3/XA9/B 0.02fF
C4796 XA1/XA3/MP3/a_216_n18# AVDD 0.07fF
C4797 XA3/XA3/MP1/a_216_n18# XA3/XA3/MP2/a_216_n18# 0.01fF
C4798 XA8/XA1/XA1/MP3/G XA8/XA1/XA1/MP3/a_216_n18# 0.07fF
C4799 XA5/XA6/MN1/a_324_n18# XA5/XA6/MN2/a_324_n18# 0.01fF
C4800 XA5/CN0 VREF 0.69fF
C4801 XB1/XA3/MP0/S AVSS 0.22fF
C4802 XA7/XA6/MP0/a_216_n18# AVDD 0.08fF
C4803 XA20/XA3/MN4/a_324_n18# XA20/XA3/N2 0.01fF
C4804 XA4/XA3/MP0/a_216_n18# AVDD 0.08fF
C4805 XA8/XA1/XA4/MN1/S AVSS 0.10fF
C4806 XA0/XA1/XA1/MP2/a_216_n18# XA0/XA1/XA1/MP1/a_216_n18# 0.01fF
C4807 XA1/XA5/MN2/a_324_n18# XA1/XA5/MN1/a_324_n18# 0.01fF
C4808 XA5/XA9/MP0/a_216_n18# XA5/XA9/A 0.14fF
C4809 SARN XB1/M5/a_324_n18# 0.01fF
C4810 XA6/XA9/A AVSS 0.31fF
C4811 XA6/EN D<3> 0.47fF
C4812 XA20/XA1/MP0/a_216_n18# XA20/XA1/MP0/a_216_334# 0.01fF
C4813 XA6/XA7/MP0/a_216_n18# AVDD 0.09fF
C4814 XA20/XA4/MP0/S XA20/XA4/MN4/a_324_n18# 0.01fF
C4815 XA0/XA4/MN0/a_324_n18# XA0/XA3/MN3/a_324_n18# 0.01fF
C4816 XA3/XA3/MP2/a_216_n18# VREF 0.03fF
C4817 XA6/XA4/MP2/a_216_n18# VREF 0.03fF
C4818 XA5/XA9/B XA5/XA9/A 0.29fF
C4819 XB2/XA3/MP2/a_216_n18# XB2/XA4/MP0/a_216_n18# 0.01fF
C4820 XA7/XA1/XA2/Y XA7/XA1/XA5/MN2/a_324_n18# 0.07fF
C4821 XA20/XA11/MN0/a_324_n18# CK_SAMPLE 0.08fF
C4822 XA1/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C4823 XA3/XA6/MP3/S AVDD 0.16fF
C4824 XA6/XA3/MP2/a_216_n18# XA6/XA3/MP3/a_216_n18# 0.01fF
C4825 XA1/XA5/MN0/a_324_n18# XA1/XA5/MN1/a_324_n18# 0.01fF
C4826 XA6/XA4/MN3/a_324_n18# XA6/XA4/A 0.15fF
C4827 XA2/XA2/A XA2/XA2/MN0/a_324_n18# 0.08fF
C4828 XB2/XA4/GNG CK_SAMPLE_BSSW 0.03fF
C4829 XA3/CP0 XA3/XA4/MN3/a_324_n18# 0.02fF
C4830 XA2/XA1/XA2/Y AVSS 0.27fF
C4831 XA20/XA3/MP5/a_216_n18# XA20/XA3/MP6/a_216_n18# 0.01fF
C4832 D<4> AVDD 1.99fF
C4833 D<5> XA1/CN0 0.02fF
C4834 XA0/XA11/MP1/S AVDD 0.19fF
C4835 XA20/XA11/MP1/a_216_n18# AVDD 0.08fF
C4836 XA8/XA3/MP0/a_216_n18# XA8/CN1 0.07fF
C4837 XA0/XA9/A XA0/XA9/MN0/a_324_n18# 0.15fF
C4838 XA6/XA9/A XA5/XA9/B 0.02fF
C4839 DONE VREF 0.14fF
C4840 XDAC2/XC128b<2>/XRES4/B AVSS 5.49fF
C4841 XA8/CN1 XA20/CNO 0.04fF
C4842 XA2/XA3/MN3/a_324_n18# XA2/XA3/MN2/a_324_n18# 0.01fF
C4843 XA0/XA3/MN1/a_324_n18# XA0/XA3/MN0/a_324_n18# 0.01fF
C4844 XDAC2/XC64b<1>/XRES1B/B SARN 1.79fF
C4845 XA8/XA2/A AVDD 1.11fF
C4846 XA20/CPO XA0/CN0 0.05fF
C4847 XA4/XA1/XA4/MN1/S XA4/XA4/A 0.02fF
C4848 XA0/XA2/MN3/a_324_n18# XA0/XA2/A 0.15fF
C4849 XA0/CP0 XA0/XA1/XA2/Y 0.02fF
C4850 XA1/XA11/MP1/S XA0/CEO 0.02fF
C4851 XA8/EN XA7/CP0 0.06fF
C4852 XDAC2/XC128b<2>/XRES8/B XDAC2/XC128a<1>/XRES8/B 0.21fF
C4853 XA6/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C4854 XA0/CP1 XA3/CN1 0.16fF
C4855 XA3/CN0 XA2/CN1 0.06fF
C4856 XA6/XA6/MP3/a_216_n18# XA6/XA7/MP0/a_216_n18# 0.01fF
C4857 XA8/XA1/XA5/MP2/a_216_n18# XA8/XA1/XA5/MP1/a_216_n18# 0.01fF
C4858 XA7/XA1/XA1/MP2/a_216_n18# XA20/CNO 0.08fF
C4859 XDAC1/XC1/XRES8/B XB1/XA3/B 0.07fF
C4860 XA6/XA9/A XA6/XA9/Y 0.04fF
C4861 SAR_IN CK_SAMPLE_BSSW 0.04fF
C4862 XA8/XA3/MP2/a_216_n18# D<0> 0.01fF
C4863 XA4/XA1/XA5/MN1/a_324_n18# XA4/XA1/XA5/MN2/a_324_n18# 0.01fF
C4864 XA4/XA1/XA2/Y D<4> 0.02fF
C4865 XA20/XA1/MP0/S AVSS 0.49fF
C4866 XDAC1/XC64a<0>/XRES16/B XDAC1/XC64a<0>/XRES8/B 1.42fF
C4867 XA2/XA3/MN0/a_324_n18# XA2/XA2/MN3/a_324_n18# 0.01fF
C4868 XA1/XA9/B XA1/XA9/A 0.29fF
C4869 XA8/XA1/XA4/MP1/S AVDD 0.15fF
C4870 EN XA0/XA1/XA5/MN2/a_324_n18# 0.08fF
C4871 XA5/XA9/A CK_SAMPLE 0.02fF
C4872 XA2/CP0 AVDD 1.49fF
C4873 XA1/XA3/MN2/a_324_n18# AVSS 0.01fF
C4874 XA5/XA12/A XA5/XA13/MP1/a_216_n18# 0.08fF
C4875 XB2/M6/a_324_n18# SAR_IN 0.01fF
C4876 XA8/CEO XA20/XA11/Y 0.02fF
C4877 XA7/XA2/MP1/a_216_n18# VREF 0.02fF
C4878 XA7/XA12/A XA7/XA12/MP0/a_216_n18# 0.07fF
C4879 XA1/XA1/XA4/MN1/a_324_n18# XA1/XA1/XA4/MN2/a_324_n18# 0.01fF
C4880 XA2/XA5/MP2/a_216_n18# VREF 0.03fF
C4881 XA8/XA6/MN1/S XA8/XA9/B 0.05fF
C4882 XDAC1/XC128b<2>/XRES1B/B XDAC1/XC128b<2>/XRES2/B 0.23fF
C4883 XA8/ENO XA8/XA1/XA5/MP1/S 0.02fF
C4884 XA3/XA5/MP2/a_216_n18# AVDD 0.07fF
C4885 XB2/XA0/MP0/a_216_n18# CK_SAMPLE_BSSW 0.07fF
C4886 XA8/XA1/XA5/MN2/S EN 0.01fF
C4887 XA6/XA1/XA5/MP1/S AVDD 0.13fF
C4888 XA7/XA9/MN1/S AVSS 0.15fF
C4889 XA6/CP0 VREF 0.77fF
C4890 XA4/CEO XA4/XA11/MP1/S 0.02fF
C4891 D<5> XA3/EN 0.08fF
C4892 XA6/XA9/A CK_SAMPLE 0.02fF
C4893 XA1/XA4/MP1/a_216_n18# AVDD 0.07fF
C4894 XA8/XA13/MP1/a_216_334# AVDD 0.17fF
C4895 XA6/XA1/XA5/MN2/S XA6/XA2/A 0.05fF
C4896 XA8/CEO XA20/XA13/MN1/a_324_n18# 0.06fF
C4897 XA8/XA1/XA1/MP3/S XA20/CPO 0.01fF
C4898 XA1/CN0 XDAC2/XC32a<0>/C1A 0.03fF
C4899 XA5/CP0 XA5/XA5/MP0/a_216_n18# 0.07fF
C4900 XDAC2/XC0/XRES16/B SARN 21.76fF
C4901 XA0/CP1 D<3> 0.02fF
C4902 XA1/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C4903 XDAC1/XC32a<0>/XRES16/B D<6> 0.04fF
C4904 XDAC2/XC64a<0>/XRES4/B XDAC2/XC32a<0>/XRES16/B 0.03fF
C4905 XA7/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C4906 XA3/XA1/XA1/MN2/a_324_n18# XA3/XA1/XA1/MN1/a_324_n18# 0.01fF
C4907 XA0/XA2/MP3/a_216_n18# AVDD 0.07fF
C4908 XA3/XA1/XA1/MN2/S XA3/EN 0.05fF
C4909 XA7/XA1/XA4/MN1/S XA7/EN 0.02fF
C4910 XA7/XA11/MP0/a_216_n18# AVDD 0.09fF
C4911 XA1/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C4912 XA3/XA11/MP1/a_216_n18# AVDD 0.08fF
C4913 XA8/XA4/MN0/a_324_n18# XA8/CN1 0.07fF
C4914 XA0/XA4/MP3/a_216_n18# VREF 0.03fF
C4915 EN XA2/XA1/XA2/Y 0.07fF
C4916 XA1/XA1/XA1/MP0/a_216_n18# XA1/XA1/XA0/MP1/a_216_n18# 0.01fF
C4917 XA1/XA11/A VREF 0.02fF
C4918 XA7/XA1/XA1/MP3/a_216_n18# AVDD 0.08fF
C4919 XA1/XA3/MN1/a_324_n18# XA1/XA3/MN2/a_324_n18# 0.01fF
C4920 XB2/XA4/MP1/a_216_334# AVDD 0.09fF
C4921 XA7/XA1/XA5/MP2/S XA7/XA2/A 0.06fF
C4922 XA0/CP0 XDAC1/XC128a<1>/XRES16/B 0.02fF
C4923 SAR_IN XB2/XA4/GNG 0.02fF
C4924 XA1/CEO XA2/XA9/Y 0.01fF
C4925 XA6/CN1 AVDD 1.31fF
C4926 XA3/XA4/MN0/a_324_n18# XA3/XA4/A 0.09fF
C4927 XA6/XA2/MN2/a_324_n18# AVSS 0.01fF
C4928 XA4/XA5/MN2/a_324_n18# XA4/XA5/MN1/a_324_n18# 0.01fF
C4929 XA6/XA1/XA4/MN0/a_324_n18# XA6/XA1/XA2/MN0/a_324_n18# 0.01fF
C4930 XDAC2/X16ab/XRES1B/B XDAC2/X16ab/XRES4/B 1.64fF
C4931 XDAC2/X16ab/XRES2/B XDAC2/X16ab/XRES8/B 1.58fF
C4932 XDAC2/XC0/XRES1A/B XDAC2/XC0/XRES4/B 0.29fF
C4933 XDAC2/XC64b<1>/XRES4/B XDAC2/XC0/XRES8/B 0.01fF
C4934 XA20/CPO XA0/XA1/XA4/MP1/S 0.02fF
C4935 AVDD XA8/XA6/MP1/S 0.13fF
C4936 XA7/XA4/MP0/a_216_n18# VREF 0.02fF
C4937 XDAC1/XC64b<1>/XRES16/B SARP 21.64fF
C4938 XA1/XA4/MP3/a_216_n18# XA1/XA5/MP0/a_216_n18# 0.01fF
C4939 XA0/XA5/MN2/a_324_n18# AVSS 0.01fF
C4940 DONE XA20/XA4/MP0/S 0.01fF
C4941 XA8/XA4/MP1/a_216_n18# XA8/CP0 0.02fF
C4942 XA1/XA1/XA2/Y XA1/XA1/XA5/MN0/a_324_n18# 0.02fF
C4943 XA3/XA6/MP1/S AVDD 0.12fF
C4944 XA5/XA12/A XA4/CEO 0.18fF
C4945 XA7/XA6/MN2/a_324_n18# XA7/XA6/MN1/a_324_n18# 0.01fF
C4946 XA0/XA4/A XA0/XA4/MP0/a_216_n18# 0.07fF
C4947 D<2> XA6/XA3/MN3/a_324_n18# 0.02fF
C4948 XA5/XA9/A XA4/XA9/A 0.01fF
C4949 XA3/XA9/MN1/a_324_n18# XA3/XA9/MN0/a_324_n18# 0.01fF
C4950 XDAC1/X16ab/XRES16/B XA3/CP0 0.02fF
C4951 XDAC1/XC32a<0>/XRES16/B SARP 21.65fF
C4952 XA5/EN D<4> 0.43fF
C4953 XA6/XA3/MP1/a_216_n18# AVDD 0.07fF
C4954 XA1/XA1/XA2/Y XA1/XA1/XA4/MN2/a_324_n18# 0.08fF
C4955 XB1/CKN XB1/XA4/MP0/a_216_n18# 0.15fF
C4956 D<6> XA20/CPO 0.05fF
C4957 XA7/XA11/MP0/a_216_n18# XA7/XA11/A 0.07fF
C4958 XA20/CNO XA6/XA1/XA1/MP3/G 0.06fF
C4959 XA0/XA4/A XA20/CPO 0.03fF
C4960 XA1/XA11/A XA1/XA11/MN0/a_324_n18# 0.09fF
C4961 XA2/XA6/MP1/a_216_n18# XA2/CN0 0.15fF
C4962 XB1/XCAPB1/XCAPB3/m3_252_308# XB1/XA3/B 0.02fF
C4963 XA20/XA2/N2 SARN 0.03fF
C4964 XB1/XA7/MN1/a_324_334# AVSS 0.08fF
C4965 XB1/XA4/MN1/a_324_n18# XB1/XA4/MN1/a_324_334# 0.01fF
C4966 XA0/XA6/MN3/a_324_n18# XA0/XA7/MN0/a_324_n18# 0.01fF
C4967 XA0/XA1/XA1/MN3/a_324_n18# XA1/EN 0.01fF
C4968 XA6/XA1/XA1/MP3/G XA6/XA1/XA1/MP3/S 0.04fF
C4969 XA5/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C4970 XA2/XA9/A XA2/XA11/A 0.01fF
C4971 D<3> XA5/XA3/MN3/a_324_n18# 0.02fF
C4972 XA0/XA1/XA4/MN2/S XA0/XA1/XA4/MP2/S 0.01fF
C4973 XA3/CEO XA3/XA9/B 0.03fF
C4974 XB2/XA4/MN1/S AVSS 0.14fF
C4975 XA3/XA11/MP1/S XA2/CEO 0.02fF
C4976 XA7/XA11/A XA7/XA11/MN1/a_324_n18# 0.07fF
C4977 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC64b<1>/XRES4/B 1.64fF
C4978 XA20/XA2/MP6/a_216_n18# XA20/XA3/CO 0.16fF
C4979 XB2/CKN XB2/XA3/MP0/S 0.54fF
C4980 XA7/XA1/XA1/MP1/a_216_n18# XA7/XA1/XA1/MP2/a_216_n18# 0.01fF
C4981 D<1> XA2/CN0 0.04fF
C4982 XA0/CP0 XA0/XA5/MN1/a_324_n18# 0.15fF
C4983 XA3/XA3/MN2/a_324_n18# AVSS 0.01fF
C4984 XA3/XA1/XA1/MN2/a_324_n18# XA3/XA1/XA1/MN3/a_324_n18# 0.01fF
C4985 XA0/XA2/A XA1/EN 0.10fF
C4986 XA8/ENO XA8/XA1/XA4/MP2/S 0.02fF
C4987 XA5/CP0 XA5/XA4/A 0.52fF
C4988 XA3/XA2/MP0/a_216_n18# XA3/XA1/XA5/MP2/a_216_n18# 0.01fF
C4989 XA4/CN0 XA4/XA2/A 0.04fF
C4990 XA7/XA4/MP2/a_216_n18# XA7/XA4/MP3/a_216_n18# 0.01fF
C4991 XA0/CP1 XA0/XA6/MP2/a_216_n18# 0.07fF
C4992 XA1/CP0 XA0/CN0 0.05fF
C4993 XDAC1/XC128a<1>/XRES1A/B AVSS 2.97fF
C4994 XA0/XA9/B VREF 0.12fF
C4995 XDAC1/XC32a<0>/XRES2/B SARP 3.05fF
C4996 XA3/XA11/MP0/a_216_n18# AVDD 0.09fF
C4997 XA20/XA9/A XA20/XA9/MN0/a_324_334# 0.08fF
C4998 XA6/CN0 XA6/XA1/XA2/Y 0.02fF
C4999 XA6/XA6/MP1/a_216_n18# D<2> 0.01fF
C5000 XA2/EN XA1/EN 1.81fF
C5001 XA2/XA4/A XA2/XA4/MP1/a_216_n18# 0.15fF
C5002 SARN XA20/XA3a/A 0.15fF
C5003 XA8/XA5/MN0/a_324_n18# XA8/XA5/MN1/a_324_n18# 0.01fF
C5004 XA3/CN0 VREF 0.69fF
C5005 XA7/XA1/XA5/MP1/S VREF 0.02fF
C5006 XA4/XA1/XA4/MP2/S EN 0.03fF
C5007 XA8/ENO XA8/XA1/XA4/MN0/a_324_n18# 0.07fF
C5008 XA7/XA1/XA5/MP0/a_216_n18# AVDD 0.08fF
C5009 XDAC1/XC32a<0>/XRES8/B XDAC1/XC64a<0>/XRES8/B 0.21fF
C5010 XA0/XA11/A XA0/XA11/MN0/a_324_n18# 0.09fF
C5011 XA2/XA2/MN2/a_324_n18# XA2/XA2/MN1/a_324_n18# 0.01fF
C5012 XA0/XA4/A XA0/XA1/XA5/MP1/S 0.02fF
C5013 DONE XA8/XA9/A 0.10fF
C5014 XDAC1/XC0/XRES8/B SARP 11.94fF
C5015 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC32a<0>/XRES4/B 1.64fF
C5016 XA20/CPO SARP 0.10fF
C5017 XA2/CN1 XA20/CNO 0.20fF
C5018 XDAC2/XC0/XRES1B/B SARN 1.94fF
C5019 XA1/XA1/XA2/MN0/a_324_n18# XA20/CPO 0.02fF
C5020 XA0/XA8/MN0/a_324_n18# XA0/XA9/MN0/a_324_n18# 0.01fF
C5021 XA1/XA1/XA2/Y XA1/XA4/A 0.19fF
C5022 XA3/XA11/MP0/a_216_n18# XA3/XA9/Y 0.08fF
C5023 XA5/XA2/MP0/a_216_n18# XA5/XA1/XA5/MP2/a_216_n18# 0.01fF
C5024 D<1> SARN 0.04fF
C5025 D<1> XA7/XA6/MP3/a_216_n18# 0.15fF
C5026 XA1/XA4/A XA1/XA1/XA5/MP1/S 0.02fF
C5027 XA4/XA1/XA4/MP0/a_216_n18# XA4/XA1/XA4/MP1/a_216_n18# 0.01fF
C5028 XA8/XA4/A AVSS 1.14fF
C5029 XA5/XA1/XA5/MN2/S AVSS 0.09fF
C5030 XA4/EN XA3/CN1 0.28fF
C5031 XA5/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C5032 XA4/XA6/MP1/a_216_n18# AVDD 0.08fF
C5033 XA1/XA2/MN0/a_324_n18# XA1/EN 0.07fF
C5034 XA5/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C5035 XA5/CP0 XA5/XA5/MP2/a_216_n18# 0.15fF
C5036 XA7/XA1/XA2/Y XA7/XA1/XA4/MN2/S 0.05fF
C5037 XA8/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C5038 XA20/XA1/MP0/S XA20/XA1/MN6/a_324_n18# 0.01fF
C5039 XA0/XA11/MN1/a_324_n18# XA0/XA11/A 0.07fF
C5040 XA0/CP0 XA0/XA6/MP0/a_216_n18# 0.08fF
C5041 XA8/XA2/A XA7/XA2/A 0.03fF
C5042 XA20/XA3/N1 SARP 0.31fF
C5043 XA7/XA6/MN3/S AVDD 0.01fF
C5044 XA7/CN1 XA7/CP0 0.03fF
C5045 XA3/XA2/MN2/a_324_n18# XA3/XA2/A 0.15fF
C5046 XA7/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C5047 XA2/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C5048 XA8/XA3/MN0/a_324_n18# XA8/XA2/A 0.07fF
C5049 XA0/XA9/Y XA0/XA11/A 0.14fF
C5050 XA2/XA5/MP0/a_216_n18# XA2/XA4/MP3/a_216_n18# 0.01fF
C5051 XA5/DONE XA5/XA9/A 0.07fF
C5052 XA2/CN0 XA3/CN1 2.47fF
C5053 XA2/XA9/A AVSS 0.31fF
C5054 XA5/XA1/XA1/MP3/G XA20/CNO 0.06fF
C5055 SAR_IP XB1/XA3/MP0/S 0.05fF
C5056 XA20/XA3/MN5/a_324_n18# XA20/XA3/MN6/a_324_n18# 0.01fF
C5057 AVDD XA1/CN0 4.39fF
C5058 XA7/XA1/XA4/MN2/a_324_n18# XA7/XA1/XA5/MN0/a_324_n18# 0.01fF
C5059 XDAC2/XC1/XRES8/B XDAC2/XC64a<0>/XRES8/B 0.21fF
C5060 XDAC1/XC128a<1>/XRES1B/B XDAC1/XC128a<1>/XRES4/B 1.64fF
C5061 XA3/EN XA2/XA1/XA4/MN0/a_324_n18# 0.07fF
C5062 XA3/CP0 XA3/XA4/A 0.57fF
C5063 XA4/XA1/XA1/MP3/G AVDD 0.63fF
C5064 XA5/XA1/XA0/MN1/a_324_n18# XA5/XA1/XA1/MN0/a_324_n18# 0.01fF
C5065 XA1/XA4/MN0/a_324_n18# XA1/CN1 0.07fF
C5066 XA7/CEO XA6/CEO 0.40fF
C5067 XA7/CN1 XA7/XA3/MP0/a_216_n18# 0.07fF
C5068 XA7/EN XA20/CPO 0.63fF
C5069 XA3/EN XA2/XA1/XA4/MP0/a_216_n18# 0.08fF
C5070 XA3/XA11/A AVSS 0.27fF
C5071 XA5/XA4/MP3/a_216_n18# AVDD 0.07fF
C5072 D<2> XA2/CN0 0.07fF
C5073 D<7> XA1/XA6/MP1/S 0.02fF
C5074 XA2/XA3/MN1/a_324_n18# XA2/XA3/MN0/a_324_n18# 0.01fF
C5075 XA7/EN XA6/XA1/XA1/MP2/a_216_n18# 0.02fF
C5076 XA4/XA3/MP3/a_216_n18# AVDD 0.07fF
C5077 XA7/XA5/MP0/a_216_n18# XA7/CP0 0.07fF
C5078 XA2/CN1 XA2/XA2/MP3/a_216_n18# 0.02fF
C5079 XA7/XA5/MP1/a_216_n18# XA7/CP0 0.15fF
C5080 XA5/CP0 VREF 0.77fF
C5081 XA20/XA2a/MN3/a_324_n18# XA20/XA3a/MN0/a_324_n18# 0.01fF
C5082 XA1/XA1/XA1/MN2/S XA1/EN 0.05fF
C5083 XA2/XA9/B XA2/XA9/A 0.29fF
C5084 XA3/XA1/XA1/MP3/G XA3/XA1/XA1/MP2/a_216_n18# 0.01fF
C5085 XA0/CP1 XA0/XA6/MP3/S 0.02fF
C5086 XA1/CP0 XA1/XA5/MP1/a_216_n18# 0.15fF
C5087 XA7/CN0 XA2/CN0 0.49fF
C5088 SARN XA3/CN1 0.19fF
C5089 XDAC2/XC32a<0>/XRES1B/B AVSS 2.96fF
C5090 XA6/XA1/XA1/MP0/a_216_n18# XA6/XA1/XA1/MP1/a_216_n18# 0.01fF
C5091 XA0/CP0 XA0/XA1/XA1/MP3/G 0.01fF
C5092 SARN XB1/XA1/MP0/G 0.01fF
C5093 XDAC1/XC128b<2>/XRES4/B XDAC1/XC128b<2>/XRES2/B 0.55fF
C5094 XA5/XA4/A XA20/CNO 0.21fF
C5095 XA3/XA3/MN2/a_324_n18# XA3/XA3/MN3/a_324_n18# 0.01fF
C5096 XA2/EN XA2/XA2/A 0.06fF
C5097 XA20/XA3/MN4/a_324_n18# XA20/XA3/N1 0.01fF
C5098 XB2/M6/a_324_n18# XB2/M7/a_324_n18# 0.01fF
C5099 XA4/XA1/XA1/MP3/G XA4/XA1/XA2/MP0/a_216_n18# 0.08fF
C5100 XDAC2/XC128a<1>/XRES8/B XDAC2/XC32a<0>/XRES4/B 0.01fF
C5101 D<7> XA20/CNO 0.06fF
C5102 XA6/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C5103 XB2/XA3/MP0/S XA0/CEIN 0.02fF
C5104 XA3/XA4/MP1/a_216_n18# XA3/XA4/A 0.15fF
C5105 XA20/XA9/Y XA20/XA2/N2 0.04fF
C5106 XA6/XA4/A D<1> 0.01fF
C5107 XA20/XA11/MN1/a_324_n18# AVSS 0.01fF
C5108 XA4/XA6/MP3/a_216_n18# XA4/XA7/MP0/a_216_n18# 0.01fF
C5109 XA20/XA13/MP1/a_216_n18# XA20/XA13/MP1/a_216_334# 0.01fF
C5110 XDAC2/XC128a<1>/XRES1B/B XDAC2/XC32a<0>/XRES1B/B 0.03fF
C5111 XDAC1/XC64a<0>/XRES16/B XDAC1/XC64a<0>/XRES1B/B 0.12fF
C5112 D<3> XA2/CN0 0.27fF
C5113 SARP XA0/CEIN 0.74fF
C5114 D<2> SARN 0.03fF
C5115 XA0/XA4/A XA0/XA1/XA5/MN1/S 0.02fF
C5116 XA0/XA2/A XA0/XA2/MP2/a_216_n18# 0.15fF
C5117 XA3/XA1/XA5/MN2/a_324_n18# XA3/EN 0.08fF
C5118 XA7/XA1/XA1/MP3/a_216_n18# XA7/XA1/XA2/MP0/a_216_n18# 0.01fF
C5119 XA4/XA1/XA5/MP1/S XA4/XA1/XA5/MP2/S 0.04fF
C5120 XA20/XA1/MN0/a_324_n18# AVSS 0.07fF
C5121 XA2/XA4/A XA1/XA4/A 0.16fF
C5122 XA2/EN XA1/XA1/XA4/MP2/S 0.02fF
C5123 XA4/XA1/XA1/MP0/a_216_n18# AVDD 0.15fF
C5124 XDAC2/XC0/XRES2/B XDAC2/XC0/XRES16/B 1.61fF
C5125 AVDD XA3/EN 5.03fF
C5126 XA4/XA1/XA4/MN2/S XA4/XA4/A 0.06fF
C5127 XA0/XA11/MP1/a_216_n18# XA0/CEIN 0.06fF
C5128 XA0/CP0 D<8> 0.14fF
C5129 XA5/XA2/A XA5/XA2/MN2/a_324_n18# 0.15fF
C5130 XA7/CN0 SARN 0.07fF
C5131 XA1/CP0 D<6> 3.42fF
C5132 XA8/XA4/A EN 0.09fF
C5133 XDAC2/XC64a<0>/XRES2/B SARN 3.05fF
C5134 XA5/XA1/XA5/MN2/S EN 0.02fF
C5135 XB1/XA5/MN1/a_324_n18# XB1/XA7/MN1/a_324_334# 0.01fF
C5136 XA20/XA2/MN1/a_324_n18# XA20/XA3/N1 0.02fF
C5137 XA1/XA1/XA2/Y XA1/XA1/XA5/MN1/S 0.05fF
C5138 XA2/XA9/A CK_SAMPLE 0.02fF
C5139 XA1/XA1/XA5/MP1/S XA1/XA1/XA5/MN1/S 0.01fF
C5140 XA20/XA9/Y XA20/XA3a/A 0.47fF
C5141 XA0/XA2/MN1/a_324_n18# D<8> 0.03fF
C5142 XA2/XA6/MN1/S AVSS 0.15fF
C5143 XA4/XA1/XA1/MN2/S XA20/CNO 0.03fF
C5144 XA7/XA9/B XA6/CEO 0.02fF
C5145 XA6/DONE AVSS 0.15fF
C5146 D<3> SARN 0.03fF
C5147 XB1/XA4/MP1/a_216_n18# XB1/XA3/B 0.01fF
C5148 XA7/XA6/MP2/a_216_n18# XA7/XA6/MP1/a_216_n18# 0.01fF
C5149 XA5/XA5/MN0/a_324_n18# XA5/XA4/MN3/a_324_n18# 0.01fF
C5150 XA5/XA6/MN1/S D<3> 0.01fF
C5151 XA20/XA9/A XA20/XA2/N2 0.08fF
C5152 XA3/CN0 XA3/XA2/A 0.04fF
C5153 XB1/M4/G XB1/M3/a_324_n18# 0.15fF
C5154 XA5/XA1/XA1/MP1/a_216_n18# XA5/XA1/XA1/MP2/a_216_n18# 0.01fF
C5155 XA6/XA1/XA1/MN1/a_324_n18# XA6/XA1/XA1/MN2/a_324_n18# 0.01fF
C5156 XDAC1/XC64a<0>/XRES8/B XDAC1/XC64a<0>/XRES2/B 1.58fF
C5157 XA4/XA1/XA2/Y XA3/EN 0.02fF
C5158 XA5/XA9/B XA5/XA6/MP3/S 0.07fF
C5159 XB2/XA3/MP0/a_216_334# XB2/XA3/MP0/a_216_n18# 0.01fF
C5160 XA1/XA6/MP1/S VREF 0.04fF
C5161 XA20/XA2/N2 XA20/XA2/MN4/a_324_n18# 0.01fF
C5162 XA5/XA3/MP0/a_216_n18# XA5/XA3/MP1/a_216_n18# 0.01fF
C5163 XB2/XCAPB1/XCAPB2/m3_324_308# XB2/XA3/B 0.02fF
C5164 AVDD XA2/XA1/XA1/MN2/S 0.05fF
C5165 XA3/XA1/XA2/MP0/a_216_n18# XA3/XA1/XA1/MP3/G 0.08fF
C5166 XDAC1/XC1/XRES4/B XDAC1/XC64a<0>/XRES16/B 0.03fF
C5167 XA2/XA9/B XA2/XA6/MN1/S 0.05fF
C5168 XA6/XA1/XA2/MN0/a_324_n18# XA7/EN 0.09fF
C5169 XA3/XA9/B XA3/XA6/MP3/S 0.07fF
C5170 XA8/XA3/MP0/a_216_n18# VREF 0.02fF
C5171 XA0/XA9/B XA0/XA9/MN1/a_324_334# 0.07fF
C5172 XA6/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C5173 XA8/ENO XA8/XA8/MN0/a_324_n18# 0.06fF
C5174 XA2/CN1 XA2/XA1/XA2/Y 0.05fF
C5175 VREF XA20/CNO 0.27fF
C5176 XA6/XA9/B XA6/XA9/MN1/a_324_n18# 0.09fF
C5177 XDAC2/XC1/XRES2/B SARN 3.05fF
C5178 XA1/CP0 SARP 0.35fF
C5179 XA20/XA9/A XA20/XA3a/A 0.18fF
C5180 XDAC2/X16ab/XRES8/B XDAC2/X16ab/XRES16/B 1.42fF
C5181 XA3/XA3/MN1/a_324_n18# D<5> 0.02fF
C5182 XA20/XA11/MN1/a_324_n18# CK_SAMPLE 0.06fF
C5183 XA0/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C5184 XA0/XA11/A XA0/CEIN 0.08fF
C5185 XA6/DONE XA6/XA9/Y 0.06fF
C5186 XA4/XA1/XA4/MN0/a_324_n18# XA4/XA1/XA2/MN0/a_324_n18# 0.01fF
C5187 XA1/XA11/MP0/a_216_n18# XA1/XA9/MP1/a_216_334# 0.01fF
C5188 XA7/XA2/MN1/a_324_n18# XA7/CN1 0.02fF
C5189 XA4/CN0 XA20/CPO 0.06fF
C5190 D<2> XA6/XA4/A 0.26fF
C5191 XA6/XA4/MN2/a_324_n18# XA6/CP0 0.01fF
C5192 XA6/XA2/MN2/a_324_n18# XA6/XA2/MN1/a_324_n18# 0.01fF
C5193 XA8/CN1 XA8/XA4/A 0.58fF
C5194 XA6/XA13/MN1/a_324_n18# XA6/XA12/A 0.07fF
C5195 XA1/XA3/MP3/a_216_n18# XA1/CN1 0.15fF
C5196 SAR_IN XB2/M7/a_324_n18# 0.01fF
C5197 XA7/XA4/MP2/a_216_n18# XA7/XA4/MP1/a_216_n18# 0.01fF
C5198 XA3/XA9/MP1/a_216_n18# AVDD 0.09fF
C5199 XDAC1/XC128a<1>/XRES4/B XDAC1/XC128b<2>/XRES16/B 0.03fF
C5200 XA6/XA13/MP1/a_216_334# AVDD 0.17fF
C5201 XA4/XA12/A XA4/XA11/MP1/S 0.06fF
C5202 XA4/XA1/XA1/MP3/G XA5/EN 0.28fF
C5203 XA0/XA1/XA4/MP2/S XA0/XA1/XA4/MP1/S 0.04fF
C5204 XB1/M4/G XB1/XA3/B 0.06fF
C5205 XA20/XA3a/MP0/a_216_n18# XA20/XA2a/MP3/a_216_n18# 0.01fF
C5206 XDAC2/XC1/XRES1B/B XDAC2/XC1/XRES2/B 0.23fF
C5207 XB1/M4/G XB1/M5/a_324_n18# 0.07fF
C5208 XA4/XA1/XA5/MN0/a_324_n18# XA4/XA1/XA4/MN2/a_324_n18# 0.01fF
C5209 XA1/XA1/XA1/MN2/a_324_n18# XA1/XA1/XA1/MN3/a_324_n18# 0.01fF
C5210 XA5/CN0 XA20/CPO 0.07fF
C5211 XA8/XA9/B XA8/XA9/MN1/a_324_n18# 0.09fF
C5212 XA5/XA11/MN1/a_324_n18# XA5/XA11/A 0.07fF
C5213 XA3/CP0 XA3/XA4/MP1/a_216_n18# 0.02fF
C5214 XA0/XA9/MN1/a_324_n18# XA0/XA9/B 0.09fF
C5215 XA1/CP0 XA1/XA5/MP3/a_216_n18# 0.15fF
C5216 XDAC2/XC128a<1>/XRES2/B XDAC2/XC128a<1>/XRES1A/B 0.25fF
C5217 XA1/XA9/B XA1/DONE 0.03fF
C5218 XA5/XA1/XA5/MP2/S EN 0.04fF
C5219 XA2/XA6/MN1/S CK_SAMPLE 0.04fF
C5220 XA1/XA9/B XA1/XA7/MN0/a_324_n18# 0.01fF
C5221 XA8/XA1/XA2/Y XA8/XA1/XA5/MN0/a_324_n18# 0.02fF
C5222 XA4/XA3/MN1/a_324_n18# XA4/XA3/MN0/a_324_n18# 0.01fF
C5223 XA2/XA9/MN1/S AVSS 0.15fF
C5224 D<1> XA7/XA3/MN1/a_324_n18# 0.02fF
C5225 D<1> D<5> 0.02fF
C5226 D<4> XA1/CN1 0.04fF
C5227 SAR_IP XB1/M8/a_324_n18# 0.01fF
C5228 XA1/EN XA0/XA1/XA1/MP2/S 0.14fF
C5229 XA0/XA4/A XA0/XA1/XA4/MP2/S 0.05fF
C5230 XA4/CP0 XA4/XA4/MN2/a_324_n18# 0.01fF
C5231 XA8/XA9/MP1/a_216_334# XA8/XA9/B 0.08fF
C5232 XA2/XA9/Y AVDD 0.58fF
C5233 XA5/XA1/XA4/MN2/S AVSS 0.06fF
C5234 XA0/XA6/MP3/a_216_n18# XA0/XA7/MP0/a_216_n18# 0.01fF
C5235 XB1/M7/a_324_n18# XA0/CEIN 0.15fF
C5236 XA8/ENO XA8/XA1/XA1/MP2/a_216_n18# 0.02fF
C5237 XA8/XA1/XA2/Y XA20/CNO 0.21fF
C5238 XA5/CN1 XA5/XA2/MN2/a_324_n18# 0.02fF
C5239 XA4/XA4/MP2/a_216_n18# XA4/XA4/MP3/a_216_n18# 0.01fF
C5240 XA2/XA2/MP3/a_216_n18# VREF 0.03fF
C5241 XDAC2/XC0/XRES1B/B XDAC2/XC0/XRES2/B 0.23fF
C5242 AVDD XB1/XA3/B 2.43fF
C5243 XA2/XA4/A XA2/XA5/MN0/a_324_n18# 0.07fF
C5244 XA5/XA9/MN1/a_324_n18# XA5/XA9/MN0/a_324_n18# 0.01fF
C5245 XA6/XA11/A AVSS 0.28fF
C5246 XA3/XA3/MP1/a_216_n18# XA3/XA3/MP0/a_216_n18# 0.01fF
C5247 XA6/XA2/MN3/a_324_n18# XA6/XA2/MN2/a_324_n18# 0.01fF
C5248 XA2/XA1/XA4/MN2/S AVSS 0.06fF
C5249 XA1/XA6/MN0/a_324_n18# AVSS 0.01fF
C5250 XB2/XA4/GNG XDAC2/XC1/XRES4/B 0.16fF
C5251 XDAC2/XC64a<0>/XRES8/B XDAC2/XC64a<0>/XRES16/B 1.42fF
C5252 XA2/XA3/MP1/a_216_n18# XA2/CN1 0.15fF
C5253 XA6/CEO AVSS 0.49fF
C5254 XA2/XA9/MN1/S XA2/XA9/B 0.02fF
C5255 XA4/XA1/XA1/MP0/a_216_n18# XA5/EN 0.01fF
C5256 XA6/XA9/A XA6/XA8/MN0/a_324_n18# 0.09fF
C5257 XDAC2/XC64b<1>/XRES1A/B XDAC2/XC64b<1>/XRES4/B 0.29fF
C5258 XDAC2/XC64b<1>/XRES2/B XDAC2/XC64b<1>/XRES1B/B 0.23fF
C5259 XA3/XA1/XA5/MN1/a_324_n18# XA20/CNO 0.07fF
C5260 XDAC2/XC128b<2>/XRES4/B XDAC2/XC128b<2>/XRES8/B 2.60fF
C5261 XDAC1/XC32a<0>/XRES8/B XDAC1/XC64a<0>/XRES1B/B 0.02fF
C5262 XA3/XA3/MP0/a_216_n18# VREF 0.02fF
C5263 XDAC1/X16ab/XRES2/B XDAC1/X16ab/XRES16/B 1.61fF
C5264 XA2/CP0 XA1/CN1 0.04fF
C5265 XA6/XA1/XA2/Y XA6/XA1/XA4/MN2/a_324_n18# 0.08fF
C5266 XA3/CEO AVSS 0.53fF
C5267 XDAC1/XC64b<1>/XRES16/B XDAC1/X16ab/XRES8/B 0.03fF
C5268 XA0/XA1/XA1/MN1/a_324_n18# XA0/XA1/XA1/MN0/a_324_n18# 0.01fF
C5269 XA6/XA1/XA2/MN0/a_324_n18# XA6/XA1/XA1/MN3/a_324_n18# 0.01fF
C5270 XA1/XA1/XA2/MP0/a_216_n18# XA1/XA1/XA1/MP3/a_216_n18# 0.01fF
C5271 XA4/XA8/MP0/a_216_n18# AVDD 0.09fF
C5272 XA4/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C5273 XA7/XA1/XA5/MN0/a_324_n18# XA20/CNO 0.09fF
C5274 XA6/XA1/XA1/MN2/S AVSS 0.30fF
C5275 XB2/XCAPB1/XCAPB3/m3_9756_132# XB2/XA3/B 0.07fF
C5276 XA6/XA2/MP0/a_216_n18# AVDD 0.08fF
C5277 XDAC1/XC128b<2>/XRES2/B AVSS 3.71fF
C5278 XA6/XA4/MP0/a_216_n18# XA6/CN1 0.08fF
C5279 XA4/XA4/A XA4/CN1 0.58fF
C5280 XA0/CP1 XA1/XA4/A 0.01fF
C5281 XB1/M1/a_324_n18# AVSS 0.02fF
C5282 XA0/XA6/MP1/S AVDD 0.12fF
C5283 XA7/XA3/MP3/a_216_n18# AVDD 0.07fF
C5284 XA1/XA9/MN1/a_324_n18# XA1/XA9/MN0/a_324_n18# 0.01fF
C5285 XA0/XA9/Y XA0/XA11/MP0/a_216_n18# 0.08fF
C5286 XA2/EN XA1/XA1/XA4/MN0/a_324_n18# 0.07fF
C5287 XA1/XA9/Y VREF 0.03fF
C5288 XA1/CN0 XDAC2/XC32a<0>/XRES16/B 0.02fF
C5289 XDAC2/XC0/XRES8/B SARP 0.02fF
C5290 XA7/XA3/MN0/a_324_n18# XA7/XA2/MN3/a_324_n18# 0.01fF
C5291 XA6/XA1/XA5/MP2/S XA7/EN 0.02fF
C5292 XA4/XA1/XA4/MN2/S XA4/XA1/XA4/MN1/S 0.04fF
C5293 XA6/EN XA4/XA4/A 0.03fF
C5294 D<5> XA3/CN1 0.87fF
C5295 XA6/XA9/Y XA6/XA11/A 0.14fF
C5296 XA1/XA4/A XA1/XA4/MN3/a_324_n18# 0.15fF
C5297 XB1/M2/a_324_n18# SAR_IP 0.02fF
C5298 XA7/XA3/MP2/a_216_n18# VREF 0.03fF
C5299 XA8/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C5300 XDAC2/XC1/XRES4/B XDAC2/XC64a<0>/XRES1A/B 0.01fF
C5301 XA5/XA9/A VREF 0.04fF
C5302 XA6/XA1/XA1/MP2/S XA6/XA1/XA1/MP3/S 0.04fF
C5303 XA0/CP1 XA0/CP0 7.62fF
C5304 XA6/XA9/Y XA6/CEO 0.01fF
C5305 XA3/XA9/B XA3/XA6/MP1/S 0.07fF
C5306 XA20/XA2/MP1/a_216_n18# XA20/XA9/Y 0.14fF
C5307 XA6/XA4/A XA8/EN 0.03fF
C5308 XA4/XA9/MP1/a_216_n18# XA4/XA9/MP0/a_216_n18# 0.01fF
C5309 XA5/XA1/XA5/MN0/a_324_n18# XA5/XA1/XA5/MN1/a_324_n18# 0.01fF
C5310 XA3/XA6/MN3/S AVDD 0.01fF
C5311 XA1/XA4/MN0/a_324_n18# AVSS 0.01fF
C5312 XA6/XA2/A XA6/EN 0.06fF
C5313 XA8/XA4/MP3/a_216_n18# XA8/XA5/MP0/a_216_n18# 0.01fF
C5314 XDAC2/XC64a<0>/XRES4/B AVSS 5.50fF
C5315 D<2> D<5> 0.02fF
C5316 XA1/XA2/A XA1/CN0 0.04fF
C5317 XA8/XA13/MP1/a_216_n18# AVDD 0.13fF
C5318 XA20/XA3/N2 XA20/CNO 0.01fF
C5319 XA1/XA1/XA5/MP2/S XA1/XA4/A 0.02fF
C5320 XDAC2/XC64b<1>/XRES2/B XDAC2/XC0/XRES16/B 0.01fF
C5321 XA6/XA9/B XA6/XA6/MP3/S 0.07fF
C5322 XA4/XA1/XA5/MN2/S AVDD 0.02fF
C5323 XA20/XA9/A XA20/XA4/MP0/a_216_334# 0.08fF
C5324 XA1/XA6/MP1/a_216_n18# XA1/XA6/MP0/a_216_n18# 0.01fF
C5325 XA3/XA2/A XA20/CNO 0.04fF
C5326 XA6/XA9/A VREF 0.04fF
C5327 VREF XA2/XA5/MP0/a_216_n18# 0.02fF
C5328 XA1/XA11/MN0/a_324_n18# XA1/XA9/Y 0.07fF
C5329 XA7/XA9/MP1/a_216_334# AVDD 0.09fF
C5330 XA6/XA5/MP2/a_216_n18# AVDD 0.07fF
C5331 XA1/XA6/MN0/a_324_n18# CK_SAMPLE 0.08fF
C5332 XA3/XA8/MP0/a_216_n18# XA4/EN 0.08fF
C5333 XA7/XA1/XA5/MN1/S XA7/XA1/XA5/MN2/S 0.04fF
C5334 AVDD XA2/XA1/XA4/MP2/S 0.11fF
C5335 XDAC1/XC1/XRES2/B XB1/XA3/B 0.05fF
C5336 XDAC1/XC1/XRES8/B XDAC1/XC1/XRES16/B 1.42fF
C5337 XDAC2/X16ab/XRES4/B AVSS 5.49fF
C5338 XA3/XA6/MN0/a_324_n18# XA3/XA6/MN1/a_324_n18# 0.01fF
C5339 D<5> D<3> 0.03fF
C5340 XA3/XA1/XA5/MN2/S XA3/CN1 0.01fF
C5341 XA8/XA11/MP1/S DONE 0.01fF
C5342 XB2/XA4/MN1/S XB2/M4/G 0.11fF
C5343 XA1/XA9/B XA1/XA6/MP3/S 0.07fF
C5344 SARN XDAC2/XC32a<0>/XRES8/B 11.94fF
C5345 XA1/XA9/B AVSS 0.61fF
C5346 XA1/CP0 XA1/XA4/MN1/a_324_n18# 0.03fF
C5347 XA8/XA1/XA1/MP3/G AVSS 0.14fF
C5348 XA1/XA9/MN1/a_324_334# XA1/XA9/B 0.07fF
C5349 XDAC1/XC64b<1>/XRES4/B XDAC1/XC0/XRES16/B 0.03fF
C5350 XA0/XA1/XA5/MP0/a_216_n18# XA0/XA1/XA4/MP2/a_216_n18# 0.01fF
C5351 XA3/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C5352 XDAC1/XC1/XRES1B/B XDAC1/XC64a<0>/XRES8/B 0.02fF
C5353 XA0/XA2/A XA0/CN0 0.03fF
C5354 XA2/XA1/XA2/MN0/a_324_n18# XA2/XA1/XA1/MN3/a_324_n18# 0.01fF
C5355 D<4> XA4/XA4/MP0/a_216_n18# 0.01fF
C5356 XA6/XA4/MN0/a_324_n18# XA6/XA3/MN3/a_324_n18# 0.01fF
C5357 XA3/XA6/MP3/a_216_n18# XA3/XA6/MP2/a_216_n18# 0.01fF
C5358 XA20/XA1/MN1/a_324_n18# SARP 0.08fF
C5359 XA0/XA9/Y XA0/XA9/B 0.15fF
C5360 XDAC2/XC128a<1>/XRES16/B XDAC2/XC128a<1>/XRES1A/B 1.60fF
C5361 AVDD XB1/XA5b/MP1/a_216_n18# 0.16fF
C5362 XA2/EN XA0/CN0 0.05fF
C5363 AVDD XA2/XA1/XA1/MP2/a_216_n18# 0.08fF
C5364 XA1/XA2/MP2/a_216_n18# VREF 0.03fF
C5365 XA20/XA3/MN0/a_324_n18# XA20/XA3a/A 0.07fF
C5366 XA3/XA9/MP0/a_216_n18# AVDD 0.09fF
C5367 XA8/XA1/XA2/Y XA8/XA1/XA4/MN1/S 0.05fF
C5368 XA8/XA1/XA5/MP2/a_216_n18# EN 0.16fF
C5369 XA1/XA9/B XA2/XA9/B 0.07fF
C5370 XA1/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C5371 XA5/XA4/MP0/a_216_n18# AVDD 0.08fF
C5372 XA8/XA8/MP0/a_216_n18# XA8/XA9/A 0.07fF
C5373 XA7/XA5/MP3/a_216_n18# VREF 0.02fF
C5374 XA20/XA3/N1 XA20/XA3a/MN0/a_324_n18# 0.01fF
C5375 XA0/XA1/XA1/MP3/a_216_n18# AVDD 0.08fF
C5376 XA3/XA1/XA5/MP2/S XA3/XA4/A 0.02fF
C5377 D<3> XA4/CP0 0.01fF
C5378 XA7/XA12/MP0/a_216_n18# AVDD 0.08fF
C5379 XB2/M3/a_324_n18# XB2/M4/G 0.15fF
C5380 XB1/M5/a_324_n18# XB1/M6/a_324_n18# 0.01fF
C5381 XA4/XA2/A XA4/XA2/MN0/a_324_n18# 0.08fF
C5382 XA20/XA3/N1 XA20/XA3a/MN3/a_324_n18# 0.01fF
C5383 XA4/XA2/A XA20/CNO 0.03fF
C5384 XA0/XA1/XA5/MP2/S XA1/EN 0.02fF
C5385 XDAC1/XC64a<0>/XRES1B/B XDAC1/XC64a<0>/XRES2/B 0.23fF
C5386 XA6/XA3/MN2/a_324_n18# XA6/XA3/MN1/a_324_n18# 0.01fF
C5387 XA5/XA8/MP0/a_216_n18# AVDD 0.09fF
C5388 XB2/XA5/MP1/a_216_n18# XB2/XA4/GNG 0.01fF
C5389 XA7/XA13/MN1/a_324_334# XA7/XA13/MN1/a_324_n18# 0.01fF
C5390 XA3/XA2/A XA3/XA3/MP0/a_216_n18# 0.08fF
C5391 XB2/XA3/MP2/a_216_n18# AVDD 0.16fF
C5392 XA4/XA8/MP0/a_216_n18# XA5/EN 0.08fF
C5393 XA7/XA1/XA5/MN2/S XA20/CNO 0.01fF
C5394 XB1/XA1/MP0/G XB1/XA4/MP1/a_216_334# 0.06fF
C5395 XA20/XA2/N2 AVDD 0.47fF
C5396 XA5/EN XA5/XA1/XA4/MN2/a_324_n18# 0.08fF
C5397 XA2/XA3/MP1/a_216_n18# VREF 0.02fF
C5398 XB2/XA4/MP0/a_216_n18# XB2/XA4/MP1/a_216_n18# 0.01fF
C5399 XA3/XA1/XA5/MN1/S XA3/XA4/A 0.02fF
C5400 XA0/XA6/MP1/a_216_n18# XA0/XA6/MP2/a_216_n18# 0.01fF
C5401 XDAC2/XC128b<2>/XRES1A/B SARN 1.50fF
C5402 XA3/CN0 XA20/CPO 0.06fF
C5403 XA7/XA11/MP1/S VREF 0.01fF
C5404 XA6/XA1/XA2/Y XA5/XA1/XA2/Y 0.02fF
C5405 XA7/XA6/MP3/a_216_n18# XA7/XA7/MP0/a_216_n18# 0.01fF
C5406 XA3/XA1/XA5/MP1/S XA3/XA4/A 0.02fF
C5407 EN XA5/XA1/XA4/MP2/S 0.03fF
C5408 XA5/XA3/MP1/a_216_n18# VREF 0.02fF
C5409 XA6/XA1/XA4/MP1/S XA6/XA1/XA4/MP2/S 0.04fF
C5410 XA6/XA1/XA2/Y XA6/XA1/XA4/MN1/S 0.05fF
C5411 D<0> XA20/XA9/Y 0.01fF
C5412 XA1/XA6/MN1/S AVSS 0.15fF
C5413 XA2/XA1/XA1/MP3/G XA2/XA1/XA2/MN0/a_324_n18# 0.06fF
C5414 XA1/XA9/B CK_SAMPLE 0.09fF
C5415 XA2/EN XA1/XA1/XA1/MN3/a_324_n18# 0.02fF
C5416 XA1/XA1/XA1/MP1/a_216_n18# EN 0.08fF
C5417 XDAC1/XC0/XRES4/B XDAC1/XC0/XRES8/B 2.60fF
C5418 XA1/XA4/MP3/a_216_n18# XA1/XA4/MP2/a_216_n18# 0.01fF
C5419 XA4/CP0 XA4/XA4/MP3/a_216_n18# 0.02fF
C5420 XA5/XA2/MN1/a_324_n18# XA5/XA2/MN2/a_324_n18# 0.01fF
C5421 XB1/XCAPB1/XCAPB1/m3_9756_132# XB1/XA4/GNG 0.02fF
C5422 XA6/XA1/XA4/MN2/S XA20/CNO 0.01fF
C5423 XA2/XA6/MP1/a_216_n18# AVDD 0.08fF
C5424 XA7/XA11/MP1/a_216_n18# XA6/CEO 0.07fF
C5425 XB2/M1/a_324_n18# AVSS 0.02fF
C5426 XA8/XA1/XA4/MP0/a_216_n18# EN 0.07fF
C5427 XA2/XA12/MN0/a_324_n18# AVSS 0.01fF
C5428 AVDD XA20/XA3a/A 3.40fF
C5429 XA2/XA1/XA1/MP1/a_216_n18# XA2/XA1/XA1/MP3/G 0.01fF
C5430 XA5/XA11/MP1/a_216_n18# AVDD 0.08fF
C5431 XA4/XA1/XA1/MN3/a_324_n18# XA4/XA1/XA2/MN0/a_324_n18# 0.01fF
C5432 XA8/XA1/XA1/MP3/G EN 0.10fF
C5433 XA5/CN0 XA5/XA6/MP2/a_216_n18# 0.08fF
C5434 XDAC1/XC32a<0>/XRES4/B XDAC1/XC128a<1>/XRES8/B 0.01fF
C5435 XB2/XA1/Y XB2/XA3/MP0/S 0.02fF
C5436 XA5/XA4/A XA5/XA1/XA5/MN2/S 0.02fF
C5437 XA3/XA9/A XA3/XA9/MN0/a_324_n18# 0.15fF
C5438 XA4/XA9/Y XA4/XA11/MN0/a_324_n18# 0.07fF
C5439 AVDD XA2/XA1/XA1/MP2/S 0.11fF
C5440 D<1> AVDD 1.99fF
C5441 XA5/XA4/MP2/a_216_n18# XA5/XA4/MP3/a_216_n18# 0.01fF
C5442 XA4/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C5443 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC64b<1>/XRES1A/B 0.01fF
C5444 XA0/XA11/MP0/a_216_n18# XA0/XA9/MP1/a_216_334# 0.01fF
C5445 XA1/CN0 XA1/CN1 1.40fF
C5446 XA7/XA1/XA1/MP3/G XA7/EN 0.09fF
C5447 XA3/XA3/MP3/a_216_n18# XA3/CN1 0.15fF
C5448 D<4> AVSS 2.25fF
C5449 XA0/XA1/XA2/Y D<8> 0.05fF
C5450 XB2/XA1/Y SARP 0.02fF
C5451 XA7/XA1/XA5/MP2/S EN 0.04fF
C5452 XA8/XA2/MP2/a_216_n18# XA8/XA2/MP3/a_216_n18# 0.01fF
C5453 XA20/XA11/MP1/a_216_n18# XA20/XA12/Y 0.01fF
C5454 XA8/XA9/A XA8/XA9/MN1/a_324_n18# 0.07fF
C5455 XA8/XA1/XA1/MN2/S XA8/XA1/XA1/MP3/G 0.08fF
C5456 XA5/XA9/MN1/a_324_n18# XA5/XA9/MN1/a_324_334# 0.01fF
C5457 XA3/XA1/XA1/MN1/a_324_n18# XA3/EN 0.07fF
C5458 XA1/XA13/MN1/a_324_n18# AVSS 0.09fF
C5459 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128a<1>/XRES4/B 2.60fF
C5460 XDAC1/XC64a<0>/XRES8/B SARP 11.94fF
C5461 XA8/XA2/A AVSS 0.30fF
C5462 XA1/XA11/A XA1/XA11/MP1/a_216_n18# 0.08fF
C5463 XA1/XA1/XA5/MN0/a_324_n18# XA1/XA1/XA5/MN1/a_324_n18# 0.01fF
C5464 XA6/XA13/MN1/a_324_n18# XA6/XA13/MN1/a_324_334# 0.01fF
C5465 XA0/XA13/MN1/a_324_334# AVSS 0.09fF
C5466 XA0/XA4/A XA0/XA2/A 0.15fF
C5467 XA2/XA8/MN0/a_324_n18# XA3/EN 0.06fF
C5468 XB1/M4/G XB1/XA1/MP0/G 0.04fF
C5469 XA1/XA2/MP2/a_216_n18# XA1/XA2/MP3/a_216_n18# 0.01fF
C5470 XA2/XA12/A XA2/XA11/MP1/S 0.06fF
C5471 XA2/EN D<6> 0.03fF
C5472 XA1/XA1/XA2/Y XA1/XA1/XA4/MN1/a_324_n18# 0.09fF
C5473 XA2/EN XA0/XA4/A 0.03fF
C5474 XA2/XA1/XA4/MP1/S XA2/XA1/XA4/MN1/S 0.01fF
C5475 D<6> XA2/XA6/MP2/a_216_n18# 0.07fF
C5476 XA4/XA11/MN0/a_324_n18# XA4/XA11/MN1/a_324_n18# 0.01fF
C5477 XA1/XA6/MN1/S CK_SAMPLE 0.05fF
C5478 XA0/XA9/B XA0/CEIN 0.02fF
C5479 XDAC2/XC64b<1>/XRES8/B XDAC2/X16ab/XRES4/B 0.01fF
C5480 XA2/CP0 AVSS 1.23fF
C5481 XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MP3/a_216_n18# 0.07fF
C5482 XA5/XA6/MP2/a_216_n18# XA5/XA6/MP3/a_216_n18# 0.01fF
C5483 XDAC1/XC128a<1>/XRES2/B SARP 3.05fF
C5484 XB1/XA3/MP0/a_216_334# XB1/XA3/B 0.02fF
C5485 XDAC2/XC64b<1>/XRES1B/B XDAC2/X16ab/XRES1B/B 0.03fF
C5486 XB2/M2/a_324_n18# XB2/M3/a_324_n18# 0.01fF
C5487 XA1/XA12/A XA1/XA11/MP1/S 0.06fF
C5488 XDAC2/XC128a<1>/XRES4/B SARN 6.32fF
C5489 XA3/XA12/MP0/a_216_n18# AVDD 0.08fF
C5490 XA5/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C5491 VREF XA8/XA5/MP1/a_216_n18# 0.02fF
C5492 XDAC1/XC32a<0>/C1A XA1/CP0 0.03fF
C5493 XA4/XA7/MP0/a_216_n18# AVDD 0.09fF
C5494 XA5/XA1/XA1/MP2/a_216_n18# XA20/CNO 0.08fF
C5495 XA7/XA6/MN0/a_324_n18# XA7/CP0 0.07fF
C5496 XA0/XA11/A XA0/XA12/A 0.07fF
C5497 XA1/XA1/XA4/MP1/S EN 0.02fF
C5498 AVDD XA3/CN1 1.39fF
C5499 XA1/XA1/XA4/MN2/S AVDD 0.02fF
C5500 XDAC1/XC128b<2>/XRES8/B XDAC1/XC128b<2>/XRES2/B 1.58fF
C5501 XA4/XA1/XA1/MN3/a_324_n18# XA20/CPO 0.08fF
C5502 AVDD XA1/XA5/MP2/a_216_n18# 0.07fF
C5503 XA8/XA6/MP2/a_216_n18# XA8/XA6/MP3/a_216_n18# 0.01fF
C5504 AVDD XB1/XA1/MP0/G 0.28fF
C5505 XA3/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C5506 XA8/XA2/MP1/a_216_n18# XA8/XA2/MP2/a_216_n18# 0.01fF
C5507 SAR_IP XB1/M1/a_324_n18# 0.01fF
C5508 XA8/XA4/A VREF 0.32fF
C5509 XA0/CP0 SARN 0.02fF
C5510 XA20/XA3/MN6/a_324_n18# SARN 0.08fF
C5511 XA8/CEO AVDD 1.52fF
C5512 D<4> CK_SAMPLE 0.10fF
C5513 XA0/XA9/B XA0/XA9/MP1/a_216_334# 0.08fF
C5514 XDAC2/XC64a<0>/XRES2/B XDAC2/XC32a<0>/XRES2/B 0.05fF
C5515 XA4/XA6/MN1/S D<4> 0.01fF
C5516 XA1/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C5517 XA5/XA4/A XA5/XA1/XA5/MP2/S 0.02fF
C5518 XA20/XA11/MP1/a_216_n18# CK_SAMPLE 0.08fF
C5519 XA0/XA3/MP1/a_216_n18# D<8> 0.15fF
C5520 D<2> AVDD 1.99fF
C5521 XA7/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C5522 XA3/XA1/XA2/Y XA3/XA4/A 0.19fF
C5523 XA6/XA2/MP1/a_216_n18# VREF 0.02fF
C5524 XA2/EN XA1/XA1/XA2/MN0/a_324_n18# 0.09fF
C5525 XA7/XA5/MN0/a_324_n18# XA7/CP0 0.09fF
C5526 XA3/XA9/B XA3/XA9/MP1/a_216_n18# 0.07fF
C5527 XA6/XA1/XA5/MN1/S XA6/XA4/A 0.02fF
C5528 XA4/XA1/XA2/Y XA3/CN1 0.03fF
C5529 XA20/XA3/MN2/a_324_n18# XA20/XA3/MN1/a_324_n18# 0.01fF
C5530 XA7/CN0 AVDD 4.70fF
C5531 XA6/XA9/B XA7/EN 0.07fF
C5532 XA5/XA11/MP0/a_216_n18# XA5/XA11/MP1/a_216_n18# 0.01fF
C5533 XA8/ENO XA20/XA9/Y 0.08fF
C5534 D<4> EN 0.07fF
C5535 XA4/XA4/A XA4/EN 0.14fF
C5536 XA6/CN0 XA6/XA5/MP1/a_216_n18# 0.02fF
C5537 XDAC1/XC32a<0>/XRES16/B XDAC1/XC64a<0>/XRES4/B 0.03fF
C5538 XA0/XA8/MP0/a_216_n18# XA0/XA7/MP0/a_216_n18# 0.01fF
C5539 XA0/XA1/XA1/MP3/G XA0/XA1/XA1/MN2/S 0.08fF
C5540 XB2/XA3/MP0/a_216_n18# CK_SAMPLE_BSSW 0.08fF
C5541 XA0/XA4/A XA0/XA4/MP2/a_216_n18# 0.15fF
C5542 XA6/CN1 AVSS 0.80fF
C5543 XDAC1/XC1/XRES8/B XDAC1/XC1/XRES1A/B 0.12fF
C5544 DONE XA8/XA9/Y 0.09fF
C5545 XA7/XA11/MN1/a_324_n18# AVSS 0.01fF
C5546 XA6/XA9/B XA5/CEO 0.02fF
C5547 XA2/XA9/A VREF 0.04fF
C5548 XA7/XA6/MN3/S XA7/XA9/B 0.09fF
C5549 XA3/XA2/MP2/a_216_n18# XA3/XA2/MP3/a_216_n18# 0.01fF
C5550 XA5/XA3/MN2/a_324_n18# XA5/XA3/MN3/a_324_n18# 0.01fF
C5551 XA6/XA1/XA1/MP3/G XA6/XA1/XA1/MN2/S 0.08fF
C5552 XA2/XA12/MN0/a_324_n18# XA2/XA12/A 0.09fF
C5553 XA20/XA3/MP2/a_216_n18# XA20/XA3a/A 0.01fF
C5554 XA3/CN0 XA1/CP0 0.17fF
C5555 XB2/XA4/GNG XB2/XCAPB1/XCAPB1/m3_252_308# 0.13fF
C5556 XA8/XA2/A EN 0.13fF
C5557 XA8/XA1/XA5/MP1/S XA8/XA1/XA5/MN1/S 0.01fF
C5558 D<3> AVDD 1.99fF
C5559 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128b<2>/XRES1B/B 0.01fF
C5560 XA20/XA3/MP5/a_216_n18# XA20/XA3a/A 0.15fF
C5561 XA4/XA1/XA5/MN0/a_324_n18# XA4/EN 0.07fF
C5562 AVDD XA20/XA4/MP0/a_216_334# 0.16fF
C5563 XA2/CP0 CK_SAMPLE 0.08fF
C5564 XA6/XA6/MP3/a_216_n18# D<2> 0.15fF
C5565 XB1/XCAPB1/XCAPB1/m3_252_308# XB1/XA4/GNG 0.13fF
C5566 XB2/XA4/MP0/a_216_n18# XB2/XA4/GNG 0.02fF
C5567 XA1/XA1/XA5/MN2/a_324_n18# XA1/XA2/MN0/a_324_n18# 0.01fF
C5568 XA4/XA1/XA4/MP2/a_216_n18# XA4/XA1/XA4/MP1/a_216_n18# 0.01fF
C5569 XA20/CPO XA20/CNO 4.11fF
C5570 XA3/XA11/A VREF 0.02fF
C5571 XA7/XA5/MN2/a_324_n18# XA7/XA5/MN1/a_324_n18# 0.01fF
C5572 XA7/XA4/MN2/a_324_n18# XA7/XA4/MN3/a_324_n18# 0.01fF
C5573 XA7/XA4/MP3/a_216_n18# XA7/XA4/A 0.15fF
C5574 XA0/CP0 XDAC1/XC1/XRES8/B 0.01fF
C5575 XA0/XA2/A XA0/XA2/MN2/a_324_n18# 0.15fF
C5576 XA6/XA1/XA1/MP2/a_216_n18# XA20/CNO 0.08fF
C5577 XA4/XA1/XA5/MN2/S XA4/XA1/XA5/MN1/S 0.04fF
C5578 XA0/XA1/XA1/MN2/S D<8> 0.01fF
C5579 XA3/XA1/XA1/MP3/G XA3/EN 0.09fF
C5580 XA8/XA1/XA2/Y XA8/XA4/A 0.19fF
C5581 XA8/XA11/MP1/a_216_n18# XA8/XA11/A 0.08fF
C5582 XA7/XA1/XA1/MN2/S AVDD 0.05fF
C5583 XA8/XA1/XA4/MP1/S EN 0.02fF
C5584 XA8/XA1/XA2/MN0/a_324_n18# XA8/XA1/XA1/MN3/a_324_n18# 0.01fF
C5585 XB1/XCAPB1/XCAPB4/m3_9828_132# XB1/XA3/B 0.21fF
C5586 XA2/CP0 EN 0.05fF
C5587 XA6/XA4/MN0/a_324_n18# XA6/XA4/A 0.09fF
C5588 XA2/CP0 XA2/XA4/MN3/a_324_n18# 0.02fF
C5589 XA8/XA1/XA0/MP1/a_216_n18# XA8/XA1/XA1/MP0/a_216_n18# 0.01fF
C5590 XA20/XA2/MP1/a_216_n18# AVDD 0.10fF
C5591 XDAC1/XC1/XRES1B/B XDAC1/XC64a<0>/XRES1B/B 0.03fF
C5592 XA2/XA9/MP0/a_216_n18# AVDD 0.09fF
C5593 XA7/XA11/MN0/a_324_n18# XA7/XA11/MN1/a_324_n18# 0.01fF
C5594 XA5/XA2/MP3/a_216_n18# AVDD 0.07fF
C5595 XA2/XA9/Y XA2/XA9/MN1/a_324_334# 0.09fF
C5596 XA20/XA3/N1 XA20/CNO 0.21fF
C5597 XA4/XA3/MP3/a_216_n18# XA4/XA4/MP0/a_216_n18# 0.01fF
C5598 XA3/CP0 XA3/XA6/MN0/a_324_n18# 0.07fF
C5599 XDAC1/XC64a<0>/XRES1A/B AVSS 2.97fF
C5600 XA8/XA1/XA4/MN2/S XA20/CNO 0.02fF
C5601 XA6/XA1/XA5/MP1/S EN 0.03fF
C5602 XA0/XA4/MP1/a_216_n18# VREF 0.02fF
C5603 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC64b<1>/XRES2/B 0.23fF
C5604 XB2/M8/a_324_n18# SAR_IN 0.01fF
C5605 XA5/XA13/MP1/a_216_n18# AVDD 0.13fF
C5606 XA4/XA4/MP3/a_216_n18# AVDD 0.07fF
C5607 XA20/XA2a/MP1/a_216_n18# XA20/XA2a/MP2/a_216_n18# 0.01fF
C5608 XB1/XA3/B XB1/XA1/Y 0.01fF
C5609 AVDD XA8/XA6/MP1/a_216_n18# 0.08fF
C5610 XA7/XA3/MN1/a_324_n18# XA7/CN1 0.16fF
C5611 XA0/XA4/MN0/a_324_n18# XA0/XA4/MN1/a_324_n18# 0.01fF
C5612 XA6/XA6/MN1/a_324_n18# XA6/XA6/MN2/a_324_n18# 0.01fF
C5613 XA5/XA1/XA5/MP2/S VREF 0.03fF
C5614 XA1/XA3/MN0/a_324_n18# XA1/XA2/MN3/a_324_n18# 0.01fF
C5615 XA4/XA9/A D<4> 0.01fF
C5616 XA8/XA2/MN3/a_324_n18# XA8/XA3/MN0/a_324_n18# 0.01fF
C5617 XA5/XA5/MP3/a_216_n18# AVDD 0.07fF
C5618 XB1/CKN XB1/XA3/B 0.29fF
C5619 XA3/XA1/XA4/MN2/S XA3/XA4/A 0.06fF
C5620 XA8/XA2/MP0/a_216_n18# XA8/XA1/XA5/MP2/a_216_n18# 0.01fF
C5621 XA1/XA12/A XA0/CEO 0.18fF
C5622 XA5/XA5/MN2/a_324_n18# AVSS 0.01fF
C5623 XA8/XA8/MN0/a_324_n18# XA8/XA7/MN0/a_324_n18# 0.01fF
C5624 XDAC1/XC128a<1>/XRES4/B XDAC1/XC128b<2>/XRES4/B 0.10fF
C5625 XA20/XA1/MN4/a_324_n18# SARP 0.16fF
C5626 XA0/XA1/XA5/MP1/S XA20/CNO 0.01fF
C5627 SARN XA20/XA4/MN6/a_324_n18# 0.07fF
C5628 XA5/XA6/MP3/S VREF 0.02fF
C5629 XDAC1/XC128a<1>/XRES1A/B XDAC1/XC128b<2>/XRES1A/B 0.03fF
C5630 XA0/CP1 XA0/XA1/XA2/Y 0.02fF
C5631 XA2/XA1/XA5/MN1/a_324_n18# XA2/XA1/XA5/MN0/a_324_n18# 0.01fF
C5632 XB2/XA4/GNG XB2/XA3/MP0/a_216_n18# 0.01fF
C5633 XA5/XA1/XA5/MN1/S XA5/XA1/XA2/Y 0.05fF
C5634 XA3/XA1/XA4/MN1/S XA20/CPO 0.04fF
C5635 XA8/XA2/A XA8/CN1 0.57fF
C5636 XA1/XA11/A XA1/XA11/MP0/a_216_n18# 0.07fF
C5637 XA4/DONE XA4/XA9/Y 0.06fF
C5638 XB2/XCAPB1/XCAPB4/m3_324_308# XB2/XA4/GNG 0.07fF
C5639 XA4/XA7/MP0/a_216_n18# XA5/EN 0.07fF
C5640 XA2/XA4/MN2/a_324_n18# XA2/XA4/MN1/a_324_n18# 0.01fF
C5641 XA3/CP0 XA3/XA1/XA2/Y 0.02fF
C5642 CK_SAMPLE XA8/XA6/MP1/S 0.01fF
C5643 XA8/EN AVDD 4.13fF
C5644 XA5/EN XA3/CN1 0.01fF
C5645 XA3/XA6/MN3/S XA3/XA9/B 0.09fF
C5646 XDAC1/XC1/XRES4/B XDAC1/XC1/XRES1B/B 1.64fF
C5647 XA3/XA6/MP1/S CK_SAMPLE 0.03fF
C5648 XA8/CN0 XA8/XA5/MP3/a_216_n18# 0.02fF
C5649 D<1> XA7/XA2/A 0.07fF
C5650 XA5/XA1/XA1/MP0/a_216_n18# XA5/XA1/XA1/MP1/a_216_n18# 0.01fF
C5651 XB1/XA4/MP1/a_216_334# XB1/XA7/MP1/a_216_n18# 0.01fF
C5652 XA1/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C5653 XA5/XA4/A XA5/XA1/XA4/MN2/S 0.06fF
C5654 SARN CK_SAMPLE_BSSW 0.01fF
C5655 XA7/XA1/XA2/MN0/a_324_n18# XA7/XA1/XA4/MN0/a_324_n18# 0.01fF
C5656 XA6/XA11/MN1/a_324_n18# XA6/XA11/A 0.07fF
C5657 XA6/CN1 EN 0.03fF
C5658 XA8/XA5/MP1/a_216_n18# XA8/CP0 0.15fF
C5659 XB2/M6/a_324_n18# SARN 0.02fF
C5660 XA4/XA4/MP2/a_216_n18# XA4/XA4/A 0.15fF
C5661 XA0/XA1/XA5/MN2/a_324_n18# XA0/XA2/MN0/a_324_n18# 0.01fF
C5662 XA0/XA6/MP2/a_216_n18# AVDD 0.09fF
C5663 XA4/XA9/MN1/a_324_n18# XA4/XA9/B 0.09fF
C5664 XA2/XA3/MP2/a_216_n18# XA2/CN1 0.15fF
C5665 XDAC2/XC128b<2>/XRES2/B XDAC2/XC128a<1>/XRES2/B 0.05fF
C5666 XB1/XCAPB1/XCAPB2/m3_324_308# XB1/XA3/B 0.02fF
C5667 XA7/XA6/MN3/S AVSS 0.13fF
C5668 XA7/XA4/MP2/a_216_n18# XA7/XA4/A 0.15fF
C5669 XA4/XA9/B XA3/XA9/A 0.02fF
C5670 XA20/XA1/MP0/a_216_n18# XA20/XA9/A 0.06fF
C5671 XA8/XA4/MN2/a_324_n18# XA8/XA4/MN1/a_324_n18# 0.01fF
C5672 XA3/XA2/MN0/a_324_n18# XA3/XA1/XA5/MN2/a_324_n18# 0.01fF
C5673 XB2/XA3/MP0/a_216_334# AVDD 0.15fF
C5674 XA8/XA4/A XA8/CP0 0.52fF
C5675 XA6/XA3/MN2/a_324_n18# XA6/CN1 0.16fF
C5676 XA7/CN0 XA5/EN 0.03fF
C5677 XA6/CN0 XA0/CN0 0.15fF
C5678 XA8/XA9/MN0/a_324_n18# XA8/XA9/MN1/a_324_n18# 0.01fF
C5679 XA4/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C5680 XA1/CN0 AVSS 1.33fF
C5681 XA2/XA6/MP3/S D<6> 0.02fF
C5682 XA5/XA11/MP1/S VREF 0.01fF
C5683 XB2/XA0/MP0/a_216_n18# XB2/XA3/MP0/a_216_n18# 0.01fF
C5684 XA20/CNO XA0/XA1/XA1/MP2/a_216_n18# 0.08fF
C5685 XB2/XA4/GNG XB2/XCAPB1/XCAPB1/m3_324_308# 0.07fF
C5686 XA4/XA1/XA1/MP3/G AVSS 0.12fF
C5687 XA4/CEO AVDD 1.41fF
C5688 XA6/XA4/MN0/a_324_n18# XA6/XA4/MN1/a_324_n18# 0.01fF
C5689 D<3> XA5/EN 0.09fF
C5690 XA0/XA1/XA1/MP3/G D<8> 0.02fF
C5691 XA1/XA2/MN1/a_324_n18# XA1/XA2/MN0/a_324_n18# 0.01fF
C5692 XA5/XA3/MP2/a_216_n18# AVDD 0.07fF
C5693 XA6/XA5/MP3/a_216_n18# VREF 0.02fF
C5694 XA6/XA1/XA4/MN0/a_324_n18# XA6/XA1/XA2/Y 0.02fF
C5695 XA0/XA1/XA4/MN1/S XA0/XA1/XA2/Y 0.05fF
C5696 XDAC1/XC64a<0>/XRES1B/B SARP 1.79fF
C5697 XA7/DONE AVDD 0.21fF
C5698 D<0> AVDD 1.85fF
C5699 XA6/XA2/A XA6/XA4/A 0.14fF
C5700 XA0/CP1 XA0/XA3/MP1/a_216_n18# 0.02fF
C5701 XDAC1/XC1/XRES16/B AVDD 0.02fF
C5702 XA8/XA1/XA4/MN1/S XA20/CPO 0.04fF
C5703 XA6/XA5/MN2/a_324_n18# XA6/XA5/MN3/a_324_n18# 0.01fF
C5704 XA5/XA2/MP0/a_216_n18# AVDD 0.08fF
C5705 XA0/CP1 XDAC1/XC128a<1>/XRES16/B 0.22fF
C5706 XA1/XA5/MP0/a_216_n18# XA1/XA5/MP1/a_216_n18# 0.01fF
C5707 XA5/XA6/MP1/a_216_n18# XA5/XA6/MP2/a_216_n18# 0.01fF
C5708 XA0/XA1/XA5/MN1/S XA20/CNO 0.01fF
C5709 XA4/XA1/XA4/MN1/S XA4/EN 0.02fF
C5710 D<6> XA2/XA1/XA1/MP3/G 0.02fF
C5711 XDAC2/XC0/XRES16/B XA1/CN1 0.01fF
C5712 XA1/CEO XA2/XA12/MP0/a_216_n18# 0.08fF
C5713 XA7/XA11/MP1/a_216_n18# XA7/XA11/MP0/a_216_n18# 0.01fF
C5714 XB2/XA4/GNG SARN 2.17fF
C5715 XA2/XA13/MN1/a_324_334# XA2/XA13/MN1/a_324_n18# 0.01fF
C5716 XA8/XA7/MP0/a_216_n18# XA8/XA8/MP0/a_216_n18# 0.01fF
C5717 D<5> XA0/CP0 0.94fF
C5718 XA20/CPO XA2/XA1/XA2/Y 0.22fF
C5719 XA2/CP0 XA2/XA4/MP3/a_216_n18# 0.02fF
C5720 XA7/XA1/XA5/MP0/a_216_n18# EN 0.16fF
C5721 XA5/XA4/A XA5/XA1/XA4/MP2/S 0.05fF
C5722 XA1/CP0 XA20/CNO 0.05fF
C5723 XA8/ENO XA8/XA1/XA5/MP2/S 0.02fF
C5724 XA7/XA1/XA1/MP2/a_216_n18# XA7/XA1/XA1/MP3/a_216_n18# 0.01fF
C5725 XDAC1/X16ab/XRES16/B SARP 21.64fF
C5726 XA0/XA9/B XA0/XA6/MN1/S 0.05fF
C5727 XA2/XA2/A XA2/XA1/XA5/MP2/S 0.06fF
C5728 XA3/EN AVSS 1.10fF
C5729 XA6/XA11/A VREF 0.02fF
C5730 XA8/XA1/XA1/MN1/a_324_n18# AVSS 0.01fF
C5731 XA8/XA1/XA4/MN1/S XA8/XA1/XA4/MN2/S 0.04fF
C5732 XDAC2/XC64b<1>/XRES1A/B XDAC2/X16ab/XRES16/B 0.04fF
C5733 XA4/XA8/MN0/a_324_n18# XA4/XA9/MN0/a_324_n18# 0.01fF
C5734 XA7/XA6/MN3/S CK_SAMPLE 0.03fF
C5735 XA7/CN0 XA7/XA2/A 0.05fF
C5736 XA7/XA4/MN1/a_324_n18# XA7/XA4/A 0.15fF
C5737 XDAC2/XC128b<2>/XRES4/B XDAC2/X16ab/XRES8/B 0.01fF
C5738 XA6/CEO VREF 0.30fF
C5739 XA6/XA3/MP0/a_216_n18# AVDD 0.08fF
C5740 XA0/XA6/MP3/S AVDD 0.16fF
C5741 XA5/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C5742 XB2/XA4/GNG XDAC2/XC1/XRES1B/B 0.03fF
C5743 XDAC2/XC32a<0>/XRES1B/B XDAC2/XC32a<0>/XRES4/B 1.64fF
C5744 XDAC2/XC32a<0>/XRES2/B XDAC2/XC32a<0>/XRES8/B 1.58fF
C5745 XA20/XA9/Y XA20/XA4/MN6/a_324_n18# 0.08fF
C5746 XA8/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C5747 XA0/CP1 XA0/XA1/XA1/MN2/S 0.02fF
C5748 SAR_IN SARN 1.04fF
C5749 XA3/XA5/MN1/a_324_n18# XA3/CN0 0.02fF
C5750 XA3/CN0 XA3/XA5/MP1/a_216_n18# 0.02fF
C5751 XDAC1/XC64b<1>/XRES4/B AVSS 5.49fF
C5752 XA1/CN0 CK_SAMPLE 0.08fF
C5753 XDAC1/XC1/XRES4/B SARP 6.32fF
C5754 XA4/XA9/B XA4/XA6/MP1/S 0.07fF
C5755 XA3/CEO VREF 0.05fF
C5756 XA20/XA1/MP0/S XA20/CPO 0.02fF
C5757 XA7/CN0 XDAC2/XC32a<0>/XRES16/B 0.02fF
C5758 XA0/XA4/MN3/a_324_n18# XA0/XA4/MN2/a_324_n18# 0.01fF
C5759 XA2/XA9/B XA3/EN 0.07fF
C5760 XA1/XA9/B D<7> 0.05fF
C5761 AVDD XB1/XA7/MP1/a_216_n18# 0.15fF
C5762 XA0/XA9/MP1/a_216_n18# XA0/XA9/A 0.08fF
C5763 XDAC2/XC64a<0>/XRES2/B XDAC2/XC32a<0>/XRES16/B 0.01fF
C5764 XDAC2/XC64a<0>/XRES1A/B SARN 1.50fF
C5765 XA5/XA6/MP0/a_216_n18# AVDD 0.08fF
C5766 XA3/XA4/MP3/a_216_n18# XA3/XA4/A 0.15fF
C5767 XA7/XA1/XA5/MP1/a_216_n18# EN 0.16fF
C5768 XA6/XA1/XA4/MP1/S AVDD 0.14fF
C5769 XA3/CP0 XA0/CN0 0.04fF
C5770 XA3/XA1/XA1/MP3/S XA4/EN 0.10fF
C5771 XA7/XA4/MP1/a_216_n18# XA7/XA4/A 0.15fF
C5772 XA4/XA6/MP1/S XA4/CN0 0.02fF
C5773 AVDD XA3/XA4/MP2/a_216_n18# 0.07fF
C5774 XDAC1/XC32a<0>/XRES4/B AVSS 5.78fF
C5775 XA2/XA9/Y XA2/XA11/A 0.14fF
C5776 D<7> XA1/XA6/MP2/a_216_n18# 0.07fF
C5777 XA20/XA3/MN2/a_324_n18# XA20/XA3/MN3/a_324_n18# 0.01fF
C5778 XA1/XA1/XA1/MP3/G AVDD 0.62fF
C5779 XA2/XA1/XA1/MN2/S AVSS 0.30fF
C5780 EN XA1/CN0 0.05fF
C5781 XA8/XA1/XA1/MP2/S XA8/XA1/XA1/MP3/G 0.04fF
C5782 XA3/XA11/MN1/a_324_n18# XA3/XA11/MN0/a_324_n18# 0.01fF
C5783 XA20/XA10/MP1/a_216_n18# XA20/XA11/Y 0.08fF
C5784 XB1/XA5/MP1/a_216_n18# XB1/XA7/MP1/a_216_334# 0.01fF
C5785 XB2/M1/a_324_n18# XB2/M4/G 0.08fF
C5786 XA4/XA1/XA1/MP3/G EN 0.10fF
C5787 D<6> XA3/XA4/A 0.01fF
C5788 XA6/CN0 XA6/XA5/MN3/a_324_n18# 0.01fF
C5789 XA20/XA1/MP0/S XA20/XA3/N1 0.01fF
C5790 XA0/CEIN XB1/XA3/MP0/S 0.02fF
C5791 XDAC2/XC1/XRES1B/B XDAC2/XC64a<0>/XRES1A/B 0.63fF
C5792 XDAC1/XC128a<1>/XRES4/B AVSS 5.49fF
C5793 D<4> XA2/CN1 0.03fF
C5794 XDAC2/XC128b<2>/XRES2/B XDAC2/XC128b<2>/XRES16/B 1.61fF
C5795 XDAC1/XC1/XRES16/B XDAC1/XC1/XRES2/B 1.61fF
C5796 XDAC1/XC64a<0>/XRES16/B XDAC1/XC64a<0>/XRES2/B 1.61fF
C5797 XA6/CN1 XA6/XA2/MN1/a_324_n18# 0.02fF
C5798 XA7/XA4/MN2/a_324_n18# AVSS 0.01fF
C5799 XA3/XA8/MP0/a_216_n18# AVDD 0.09fF
C5800 XA8/XA2/MP0/a_216_n18# XA8/XA2/A 0.08fF
C5801 XA3/EN CK_SAMPLE 0.09fF
C5802 XA7/XA2/MP0/a_216_n18# AVDD 0.08fF
C5803 XA0/XA9/B XA0/XA12/A 0.01fF
C5804 XA2/XA3/MP2/a_216_n18# VREF 0.03fF
C5805 XA3/XA1/XA4/MP2/S XA3/XA4/A 0.05fF
C5806 XA0/XA1/XA2/MP0/a_216_n18# XA0/XA1/XA1/MP3/a_216_n18# 0.01fF
C5807 XA6/EN XA6/XA1/XA1/MN0/a_324_n18# 0.08fF
C5808 XA2/XA4/MP1/a_216_n18# AVDD 0.07fF
C5809 XA8/EN XA7/XA1/XA2/MP0/a_216_n18# 0.08fF
C5810 XA3/XA1/XA5/MP2/S XA3/XA1/XA5/MP1/S 0.04fF
C5811 XA8/XA12/A XA8/XA12/MN0/a_324_n18# 0.09fF
C5812 XA7/XA9/MP1/a_216_334# XA7/XA9/B 0.08fF
C5813 XA7/XA6/MP3/S AVDD 0.16fF
C5814 XA7/XA7/MP0/a_216_n18# AVDD 0.09fF
C5815 XB1/XCAPB1/XCAPB4/m3_324_308# XB1/XA3/B 0.02fF
C5816 XA4/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C5817 XA1/XA6/MN1/S D<7> 0.01fF
C5818 XA3/XA5/MP3/a_216_n18# XA3/CP0 0.15fF
C5819 XB2/M8/a_324_n18# XB2/M7/a_324_n18# 0.01fF
C5820 XA2/CP0 XA2/CN1 0.13fF
C5821 EN XA3/EN 1.04fF
C5822 D<1> XA1/CN1 0.05fF
C5823 CK_SAMPLE_BSSW XB1/XA5b/MN1/a_324_n18# 0.01fF
C5824 XDAC1/XC32a<0>/XRES16/B XDAC1/XC128a<1>/XRES1A/B 0.04fF
C5825 XA7/CN1 AVDD 1.31fF
C5826 XA8/EN XA7/XA2/A 0.10fF
C5827 XA1/XA9/B VREF 0.12fF
C5828 XA3/XA1/XA1/MP0/a_216_n18# AVDD 0.14fF
C5829 XA4/XA9/Y XA4/XA9/MP1/a_216_334# 0.07fF
C5830 XA8/ENO AVDD 5.42fF
C5831 XA8/XA1/XA1/MP3/G XA8/XA1/XA1/MN3/a_324_n18# 0.08fF
C5832 D<7> XA1/XA3/MP3/a_216_n18# 0.02fF
C5833 XA7/XA1/XA1/MN1/a_324_n18# XA7/EN 0.07fF
C5834 XA3/XA1/XA5/MN1/S XA3/XA1/XA5/MP1/S 0.01fF
C5835 XA2/XA9/Y AVSS 0.22fF
C5836 XA6/CN0 SARP 0.02fF
C5837 XA4/CP0 XA4/XA4/A 0.52fF
C5838 VREF XA2/XA11/MP1/S 0.01fF
C5839 XA20/XA2/MN3/a_324_n18# SARP 0.15fF
C5840 XA0/XA9/MP1/a_216_n18# AVDD 0.09fF
C5841 XB1/XA3/B AVSS 5.15fF
C5842 XA7/XA1/XA5/MP2/S VREF 0.03fF
C5843 XA6/XA2/MN3/a_324_n18# XA6/CN1 0.03fF
C5844 XA7/XA9/Y XA7/XA9/MN1/S 0.12fF
C5845 XA1/XA1/XA5/MP2/S XA1/XA1/XA5/MP1/S 0.04fF
C5846 XDAC1/XC64b<1>/XRES8/B XDAC1/XC0/XRES1A/B 0.03fF
C5847 XDAC1/XC64b<1>/XRES1B/B XDAC1/XC0/XRES1B/B 0.03fF
C5848 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC64a<0>/XRES16/B 0.12fF
C5849 XA0/XA1/XA5/MN2/S D<8> 0.01fF
C5850 D<6> XA2/XA3/MN3/a_324_n18# 0.02fF
C5851 XA0/XA4/A XA0/XA1/XA5/MP2/S 0.02fF
C5852 XA1/EN XA0/XA1/XA1/MP1/a_216_n18# 0.01fF
C5853 XA6/XA4/MP0/a_216_n18# D<2> 0.01fF
C5854 XA2/XA9/MN1/a_324_n18# XA2/XA9/A 0.07fF
C5855 XA0/CP1 XA0/XA1/XA1/MP3/G 0.01fF
C5856 XB1/CKN XB1/XA3/MN1/a_324_n18# 0.15fF
C5857 XA5/XA4/A D<4> 0.01fF
C5858 XA1/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C5859 XA7/XA5/MP1/a_216_n18# AVDD 0.07fF
C5860 XA7/XA5/MP0/a_216_n18# AVDD 0.08fF
C5861 XA3/CP0 XA3/XA4/MP3/a_216_n18# 0.02fF
C5862 XA4/XA9/B XA4/XA9/Y 0.15fF
C5863 XA6/EN XA4/CN1 0.03fF
C5864 D<7> D<4> 0.06fF
C5865 XA2/XA9/B XA2/XA9/Y 0.15fF
C5866 XA4/XA5/MP3/a_216_n18# XA4/XA6/MP0/a_216_n18# 0.01fF
C5867 XA8/XA9/MP1/a_216_334# XA8/XA11/MP0/a_216_n18# 0.01fF
C5868 XA20/CNO XA2/XA1/XA5/MP1/S 0.01fF
C5869 XA2/XA7/MP0/a_216_n18# XA3/EN 0.07fF
C5870 XA2/XA6/MN1/a_324_n18# XA2/XA6/MN0/a_324_n18# 0.01fF
C5871 XA6/XA1/XA5/MN1/S AVDD 0.02fF
C5872 XDAC2/XC64b<1>/XRES1B/B AVSS 2.95fF
C5873 XDAC1/XC128b<2>/XRES2/B XDAC1/XC128b<2>/XRES1A/B 0.25fF
C5874 XA6/XA1/XA5/MN2/S XA6/XA4/A 0.02fF
C5875 AVDD XA2/XA9/MP1/a_216_334# 0.09fF
C5876 XA4/XA6/MP2/a_216_n18# D<4> 0.07fF
C5877 D<6> XA3/CP0 0.06fF
C5878 XA3/XA4/MN2/a_324_n18# XA3/XA4/MN3/a_324_n18# 0.01fF
C5879 XB1/XA1/MP0/G XB1/XA1/Y 0.13fF
C5880 AVDD XA8/CN0 1.05fF
C5881 XDAC2/X16ab/XRES1A/B SARN 1.50fF
C5882 XA0/CP1 D<8> 1.60fF
C5883 XB2/M2/a_324_n18# XB2/M1/a_324_n18# 0.01fF
C5884 CK_SAMPLE_BSSW XB1/XA0/MN0/a_324_n18# 0.08fF
C5885 XB1/CKN XB1/XA1/MP0/G 0.03fF
C5886 AVDD XA2/XA1/XA4/MP1/S 0.14fF
C5887 XDAC2/XC128b<2>/XRES16/B XDAC2/XC128a<1>/XRES2/B 0.01fF
C5888 XA3/CN1 XA1/CN1 0.29fF
C5889 XA6/CN0 XA7/EN 0.15fF
C5890 XA1/XA5/MN2/a_324_n18# AVSS 0.01fF
C5891 XB2/M4/G XB2/XA4/MP1/a_216_334# 0.08fF
C5892 XA1/XA2/MP1/a_216_n18# XA1/XA2/MP0/a_216_n18# 0.01fF
C5893 XA4/XA11/MP1/a_216_n18# XA4/XA11/MP0/a_216_n18# 0.01fF
C5894 XA0/XA4/MP2/a_216_n18# XA0/XA4/MP3/a_216_n18# 0.01fF
C5895 XA0/CP0 XA0/XA5/MP1/a_216_n18# 0.15fF
C5896 XA4/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C5897 XDAC2/XC1/XRES1A/B XDAC2/XC1/XRES2/B 0.25fF
C5898 XA4/XA1/XA1/MN2/S D<4> 0.02fF
C5899 XA5/XA1/XA1/MN1/a_324_n18# XA20/CNO 0.07fF
C5900 XA2/CP0 D<7> 0.05fF
C5901 XA4/XA9/A XA4/XA9/MN0/a_324_n18# 0.15fF
C5902 XA3/XA6/MN3/a_324_n18# CK_SAMPLE 0.15fF
C5903 XB2/M8/a_324_n18# XB2/M8/a_324_334# 0.01fF
C5904 XA3/XA1/XA1/MP1/a_216_n18# XA3/XA1/XA1/MP2/a_216_n18# 0.01fF
C5905 XDAC2/XC128a<1>/XRES2/B XDAC2/XC128a<1>/XRES16/B 1.61fF
C5906 XA5/XA1/XA4/MN1/S XA5/XA1/XA2/Y 0.05fF
C5907 XA3/XA6/MN3/S AVSS 0.13fF
C5908 XA0/XA11/A XA0/CEO 0.02fF
C5909 XA4/XA5/MN1/a_324_n18# XA4/CP0 0.15fF
C5910 XA1/XA3/MP3/a_216_n18# VREF 0.03fF
C5911 XA0/XA1/XA5/MN0/a_324_n18# XA0/XA1/XA5/MN1/a_324_n18# 0.01fF
C5912 D<2> XA1/CN1 0.04fF
C5913 XA8/XA4/A XA20/CPO 0.04fF
C5914 XA20/XA1/MP0/a_216_n18# AVDD 0.15fF
C5915 XA4/XA9/MP1/a_216_n18# XA4/XA9/MP1/a_216_334# 0.01fF
C5916 XA8/ENO XA8/XA1/XA1/MP3/a_216_n18# 0.02fF
C5917 XA7/XA6/MP0/a_216_n18# VREF 0.01fF
C5918 XA6/XA1/XA2/Y XA7/EN 0.10fF
C5919 XA4/XA3/MP0/a_216_n18# VREF 0.02fF
C5920 XA5/XA4/MN3/a_324_n18# XA5/XA4/MN2/a_324_n18# 0.01fF
C5921 XA4/XA6/MN2/a_324_n18# XA4/XA6/MN1/a_324_n18# 0.01fF
C5922 XA0/CP0 XA0/XA5/MN3/a_324_n18# 0.15fF
C5923 XA20/XA3a/A XA20/XA3a/MP3/a_216_n18# 0.16fF
C5924 XA4/XA1/XA5/MN2/S AVSS 0.09fF
C5925 XA1/XA4/A AVDD 1.42fF
C5926 XA8/XA4/MN3/a_324_n18# XA8/XA4/A 0.15fF
C5927 XA7/CN0 XA1/CN1 0.05fF
C5928 XB1/XA3/MN0/a_324_n18# XB1/XA3/MN1/a_324_n18# 0.01fF
C5929 XA6/XA3/MP2/a_216_n18# AVDD 0.07fF
C5930 XA3/XA6/MP3/S VREF 0.02fF
C5931 AVDD XA20/XA3a/MP1/a_216_n18# 0.08fF
C5932 XA3/CP0 SARP 0.05fF
C5933 XA1/XA4/A XA1/XA1/XA5/MN2/S 0.02fF
C5934 XA3/XA6/MN3/a_324_n18# XA3/XA7/MN0/a_324_n18# 0.01fF
C5935 XDAC2/XC0/XRES4/B XDAC2/XC0/XRES8/B 2.60fF
C5936 XDAC2/XC0/XRES16/B AVSS 15.94fF
C5937 XA7/XA1/XA1/MP3/G XA20/CNO 0.06fF
C5938 D<4> VREF 1.75fF
C5939 VREF XA0/XA11/MP1/S 0.01fF
C5940 D<3> XA1/CN1 0.04fF
C5941 XB1/CKN XB1/XA4/MN0/a_324_n18# 0.09fF
C5942 XA0/CP0 AVDD 1.49fF
C5943 XA8/XA1/XA4/MN2/S XA8/XA4/A 0.06fF
C5944 XA5/XA6/MN3/S AVDD 0.01fF
C5945 XA4/XA9/MP1/a_216_n18# XA4/XA9/B 0.07fF
C5946 XA0/CEIN XB1/M8/a_324_n18# 0.15fF
C5947 XA4/XA6/MP0/a_216_n18# XA4/CN0 0.08fF
C5948 D<1> XA7/XA9/B 0.05fF
C5949 XA1/XA6/MP0/a_216_n18# XA1/XA5/MP3/a_216_n18# 0.01fF
C5950 XA5/XA6/MP1/S AVDD 0.12fF
C5951 XA6/XA6/MN1/S AVDD 0.01fF
C5952 XA5/XA2/MP2/a_216_n18# AVDD 0.07fF
C5953 XA8/XA2/A VREF 0.33fF
C5954 XDAC2/XC64a<0>/XRES4/B XDAC2/XC32a<0>/XRES4/B 0.10fF
C5955 XDAC1/XC64b<1>/XRES2/B XDAC1/XC0/XRES16/B 0.01fF
C5956 XA6/XA4/A XA6/XA4/MP1/a_216_n18# 0.15fF
C5957 XA20/CNO XA2/XA1/XA1/MN1/a_324_n18# 0.07fF
C5958 XA0/XA6/MP1/S CK_SAMPLE 0.03fF
C5959 XA2/XA4/MN0/a_324_n18# XA2/XA3/MN3/a_324_n18# 0.01fF
C5960 XB2/XA4/MN1/S XA0/CEIN 0.01fF
C5961 XA0/CP0 XDAC1/XC128b<2>/XRES16/B 0.18fF
C5962 XA6/CN1 XA5/XA4/A 0.04fF
C5963 XB2/XA4/MP1/a_216_n18# AVDD 0.09fF
C5964 XA20/CNO XA2/XA1/XA5/MN1/S 0.01fF
C5965 XA3/XA1/XA1/MP3/G XA3/CN1 0.02fF
C5966 XA3/XA1/XA5/MN1/S XA3/XA1/XA2/Y 0.05fF
C5967 XB2/XA3/MN1/a_324_n18# AVSS 0.01fF
C5968 XA5/XA9/MN0/a_324_n18# XA5/XA9/B 0.01fF
C5969 XA2/XA9/Y XA2/XA12/A 0.02fF
C5970 XA3/XA11/MN0/a_324_n18# XA3/XA9/MN1/a_324_334# 0.01fF
C5971 XA5/XA1/XA5/MN1/S XA5/XA1/XA5/MP1/S 0.01fF
C5972 XA20/XA2/MP6/a_216_n18# XA20/XA2/MP6/a_216_334# 0.01fF
C5973 XA1/XA11/MP0/a_216_n18# XA1/XA9/Y 0.08fF
C5974 XB2/M7/a_324_n18# SARN 0.01fF
C5975 XB1/XA5b/MP1/a_216_n18# AVSS 0.02fF
C5976 XA4/XA1/XA1/MN2/a_324_n18# XA4/XA1/XA1/MN3/a_324_n18# 0.01fF
C5977 XDAC2/XC64a<0>/XRES8/B XDAC2/XC64a<0>/XRES4/B 2.60fF
C5978 XA8/XA1/XA2/MN0/a_324_n18# XA20/CPO 0.01fF
C5979 XA6/XA2/MP0/a_216_n18# EN 0.08fF
C5980 XDAC2/XC32a<0>/XRES8/B XDAC2/XC32a<0>/XRES16/B 1.42fF
C5981 XA8/XA1/XA1/MP0/a_216_n18# AVDD 0.15fF
C5982 XA8/XA6/MP1/S XA8/XA9/B 0.07fF
C5983 XA0/XA7/MN0/a_324_n18# XA1/EN 0.08fF
C5984 XA4/XA1/XA4/MN2/S XA4/EN 0.02fF
C5985 XA0/XA4/MP1/a_216_n18# XA0/XA4/MP0/a_216_n18# 0.01fF
C5986 XA2/XA4/A XA2/XA1/XA5/MN2/S 0.02fF
C5987 XA2/CP0 VREF 0.83fF
C5988 XA4/XA12/A AVDD 0.44fF
C5989 XA0/XA3/MN3/a_324_n18# D<8> 0.15fF
C5990 XA3/XA6/MN3/S CK_SAMPLE 0.03fF
C5991 XA4/XA6/MN1/a_324_n18# XA4/XA6/MN0/a_324_n18# 0.01fF
C5992 XA2/XA1/XA2/Y XA2/XA1/XA4/MN2/a_324_n18# 0.08fF
C5993 XA0/XA4/MN0/a_324_n18# AVSS 0.01fF
C5994 XA1/XA1/XA1/MP3/S XA1/XA1/XA1/MP2/S 0.04fF
C5995 XA8/XA5/MP0/a_216_n18# AVDD 0.08fF
C5996 XDAC2/XC128a<1>/XRES8/B XDAC2/XC128a<1>/XRES1A/B 0.12fF
C5997 XB2/XA3/MP2/a_216_n18# XB2/XA3/B 0.02fF
C5998 XA3/XA5/MP2/a_216_n18# VREF 0.03fF
C5999 XDAC1/XC1/XRES1B/B XDAC1/XC64a<0>/XRES16/B 0.05fF
C6000 XA6/XA1/XA5/MP1/S VREF 0.02fF
C6001 XA1/XA4/MP1/a_216_n18# VREF 0.02fF
C6002 AVDD XA2/XA12/MP0/a_216_n18# 0.08fF
C6003 XA1/EN XA0/CN0 0.27fF
C6004 XA20/XA2/MN6/a_324_n18# XA20/XA2/MN6/a_324_334# 0.01fF
C6005 XA7/XA2/MP0/a_216_n18# XA7/XA2/A 0.08fF
C6006 XA5/XA5/MP0/a_216_n18# XA5/XA4/MP3/a_216_n18# 0.01fF
C6007 XA5/XA1/XA2/Y XA5/XA1/XA4/MP1/S 0.01fF
C6008 XA4/XA9/MN1/a_324_n18# XA4/XA9/MN1/a_324_334# 0.01fF
C6009 XA6/XA8/MP0/a_216_n18# AVDD 0.09fF
C6010 XA1/XA1/XA2/MP0/a_216_n18# XA2/EN 0.08fF
C6011 XA20/XA2/N2 AVSS 0.22fF
C6012 XA8/XA9/MP1/a_216_334# XA8/XA9/Y 0.07fF
C6013 XA6/CN0 XA4/CN0 0.66fF
C6014 XA20/XA2/MN5/a_324_n18# SARP 0.15fF
C6015 XA8/XA1/XA2/Y XA8/XA2/A 0.01fF
C6016 XA2/CN1 XA1/CN0 2.92fF
C6017 XDAC2/XC64b<1>/XRES16/B D<8> 0.05fF
C6018 D<5> XA3/XA6/MP2/a_216_n18# 0.07fF
C6019 XA7/XA1/XA2/Y AVDD 0.33fF
C6020 XA20/XA9/A XA20/XA1/MP0/a_216_334# 0.08fF
C6021 XDAC1/XC1/XRES2/B XDAC1/XC1/XRES1A/B 0.25fF
C6022 XA5/XA9/MP0/a_216_n18# XA5/XA8/MP0/a_216_n18# 0.01fF
C6023 XA4/XA1/XA5/MN2/S EN 0.02fF
C6024 XB1/M4/G XB1/XA4/MN1/S 0.11fF
C6025 XA6/EN XA5/XA1/XA1/MN3/a_324_n18# 0.02fF
C6026 XA20/XA3/MP1/a_216_n18# XA20/XA9/Y 0.14fF
C6027 XA4/XA4/MN2/a_324_n18# AVSS 0.01fF
C6028 XA0/XA2/MP3/a_216_n18# VREF 0.03fF
C6029 XA6/CN0 XA5/CN0 3.89fF
C6030 XA5/XA2/A XA5/XA1/XA2/Y 0.01fF
C6031 XA4/XA4/A AVDD 1.42fF
C6032 XA3/XA1/XA1/MP3/a_216_n18# XA3/XA1/XA1/MP2/a_216_n18# 0.01fF
C6033 XA6/XA9/A XA7/XA9/A 0.01fF
C6034 XB1/M4/G CK_SAMPLE_BSSW 0.02fF
C6035 XA7/CN1 XA7/XA2/A 0.57fF
C6036 SAR_IN XB2/M4/a_324_n18# 0.02fF
C6037 XA5/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C6038 XA5/CN1 XA5/XA3/MP3/a_216_n18# 0.15fF
C6039 XB2/XCAPB1/XCAPB0/m3_324_308# XB2/XA3/B 0.02fF
C6040 XA4/XA1/XA1/MN2/a_324_n18# XA20/CNO 0.07fF
C6041 XA4/XA1/XA1/MP2/a_216_n18# XA5/EN 0.02fF
C6042 XA7/XA1/XA4/MP1/S XA7/XA1/XA4/MP2/S 0.04fF
C6043 XA5/XA2/A XA5/XA2/MP1/a_216_n18# 0.15fF
C6044 XA4/XA5/MN2/a_324_n18# XA4/CP0 0.15fF
C6045 XA6/XA5/MN2/a_324_n18# XA6/CP0 0.15fF
C6046 XA6/XA2/A XA6/XA2/MP2/a_216_n18# 0.15fF
C6047 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC0/XRES1A/B 0.63fF
C6048 XA6/XA6/MN0/a_324_n18# XA6/XA5/MN3/a_324_n18# 0.01fF
C6049 XDAC2/XC64b<1>/XRES1B/B XDAC2/XC64b<1>/XRES8/B 0.12fF
C6050 XA1/XA1/XA5/MN1/S AVDD 0.02fF
C6051 XDAC1/XC128a<1>/XRES4/B XDAC1/XC128b<2>/XRES8/B 0.01fF
C6052 XA6/XA1/XA4/MP0/a_216_n18# XA7/EN 0.08fF
C6053 EN XA2/XA1/XA4/MP2/S 0.03fF
C6054 XA8/XA1/XA4/MP1/S XA8/XA1/XA2/Y 0.01fF
C6055 XA4/XA8/MP0/a_216_n18# XA4/XA9/A 0.07fF
C6056 XA5/XA6/MN1/a_324_n18# XA5/XA6/MN0/a_324_n18# 0.01fF
C6057 XA0/XA1/XA2/MN0/a_324_n18# XA0/XA1/XA4/MN0/a_324_n18# 0.01fF
C6058 XA4/XA1/XA4/MP1/S XA4/XA1/XA4/MP2/S 0.04fF
C6059 XDAC1/X16ab/XRES8/B XDAC1/X16ab/XRES16/B 1.42fF
C6060 XA6/XA13/MN1/a_324_n18# AVSS 0.09fF
C6061 XA20/XA3a/A AVSS 0.27fF
C6062 XA8/XA12/MP0/a_216_n18# XA8/XA13/MP1/a_216_n18# 0.01fF
C6063 XA6/XA2/A AVDD 1.07fF
C6064 XB2/XA4/MP1/a_216_334# XB2/XA1/MP0/G 0.06fF
C6065 SAR_IP XB1/M3/a_324_n18# 0.02fF
C6066 XDAC2/XC128b<2>/XRES16/B XDAC2/XC128a<1>/XRES16/B 0.41fF
C6067 XDAC1/XC64a<0>/XRES8/B XDAC1/XC64a<0>/XRES4/B 2.60fF
C6068 XA7/CN0 XA7/XA9/B 0.07fF
C6069 XA6/CN1 VREF 0.76fF
C6070 XA4/XA11/A AVDD 0.45fF
C6071 XA4/XA1/XA4/MN2/a_324_n18# XA4/EN 0.08fF
C6072 XDAC2/XC128b<2>/XRES1B/B XDAC2/X16ab/XRES1A/B 0.63fF
C6073 XDAC2/XC128b<2>/XRES2/B XDAC2/X16ab/XRES2/B 0.05fF
C6074 XA1/XA1/XA5/MN2/S XA1/XA1/XA5/MN1/S 0.04fF
C6075 XA3/XA1/XA4/MN2/a_324_n18# XA3/XA1/XA2/Y 0.08fF
C6076 VREF XA8/XA6/MP1/S 0.04fF
C6077 XDAC2/XC0/XRES1B/B AVSS 2.91fF
C6078 AVDD XB1/XA4/MN1/S 0.01fF
C6079 XDAC2/XC1/XRES4/B SARN 6.32fF
C6080 XA4/XA1/XA2/Y XA4/XA4/A 0.19fF
C6081 D<1> AVSS 3.25fF
C6082 XA3/XA6/MP1/S VREF 0.04fF
C6083 D<2> XA6/XA6/MP2/a_216_n18# 0.07fF
C6084 XA20/XA3a/A XA20/XA3a/MP2/a_216_n18# 0.16fF
C6085 XA20/XA1/MP5_DMY/a_216_n18# AVDD 0.24fF
C6086 XA5/XA4/MN0/a_324_n18# XA5/CN1 0.07fF
C6087 XA20/XA3/MN5/a_324_n18# SARN 0.16fF
C6088 XA20/XA2a/MP3/a_216_n18# XA20/XA3/CO 0.16fF
C6089 AVDD CK_SAMPLE_BSSW 8.81fF
C6090 XA5/XA7/MN0/a_324_n18# XA6/EN 0.08fF
C6091 XA8/EN XA7/XA1/XA1/MN2/a_324_n18# 0.01fF
C6092 XA3/XA6/MN2/a_324_n18# AVSS 0.01fF
C6093 XA7/XA1/XA5/MP2/S XA7/XA1/XA5/MN2/S 0.01fF
C6094 XA0/XA2/A XA20/CNO 0.03fF
C6095 XA1/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C6096 XA4/XA1/XA2/Y XA4/XA1/XA5/MN0/a_324_n18# 0.02fF
C6097 XA2/CN1 XA3/EN 0.12fF
C6098 XA6/XA3/MP1/a_216_n18# VREF 0.02fF
C6099 XA20/XA3/MP4/a_216_n18# XA20/XA3/CO 0.02fF
C6100 XA8/XA6/MP0/a_216_n18# XA8/XA6/MP1/a_216_n18# 0.01fF
C6101 XA4/XA6/MP2/a_216_n18# XA4/XA6/MP1/a_216_n18# 0.01fF
C6102 XA7/XA1/XA1/MP1/a_216_n18# XA7/XA1/XA1/MP3/G 0.01fF
C6103 XA3/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C6104 XA4/XA12/MP0/a_216_n18# XA4/XA12/A 0.07fF
C6105 XA2/XA4/A XA4/EN 0.03fF
C6106 XA1/XA1/XA4/MP0/a_216_n18# EN 0.07fF
C6107 XA0/XA2/MN3/a_324_n18# XA0/XA2/MN2/a_324_n18# 0.01fF
C6108 XA2/EN XA20/CNO 1.02fF
C6109 XDAC2/XC1/XRES1B/B XDAC2/XC1/XRES4/B 1.64fF
C6110 XA8/XA11/A AVDD 0.45fF
C6111 SARP XA20/XA3/CO 0.05fF
C6112 XA1/XA1/XA2/Y XA1/XA1/XA5/MN1/a_324_n18# 0.08fF
C6113 XA5/XA1/XA5/MN2/a_324_n18# XA5/XA1/XA2/Y 0.07fF
C6114 XA20/XA1/MP0/S XA20/XA1/MN1/a_324_n18# 0.01fF
C6115 XDAC2/XC0/XRES1A/B XDAC2/XC0/XRES16/B 1.60fF
C6116 XA2/CN0 D<8> 0.11fF
C6117 XA3/XA12/A AVDD 0.44fF
C6118 XDAC2/XC64b<1>/XRES8/B XDAC2/XC0/XRES16/B 0.03fF
C6119 XA20/CPO XA2/XA1/XA4/MN1/a_324_n18# 0.08fF
C6120 D<7> XA1/CN0 0.49fF
C6121 XA2/CN0 XA2/XA5/MP1/a_216_n18# 0.02fF
C6122 AVDD XA2/XA1/XA1/MP3/a_216_n18# 0.08fF
C6123 XA8/XA1/XA1/MN0/a_324_n18# XA8/XA1/XA1/MN1/a_324_n18# 0.01fF
C6124 XB1/XA3/MN1/a_324_n18# AVSS 0.01fF
C6125 SAR_IP XB1/XA3/B 0.23fF
C6126 SAR_IP XB1/M5/a_324_n18# 0.02fF
C6127 XA0/XA1/XA4/MP1/S XA1/EN 0.02fF
C6128 XA3/XA1/XA2/MP0/a_216_n18# XA3/XA1/XA1/MP3/a_216_n18# 0.01fF
C6129 XA4/CN0 XA3/CP0 0.04fF
C6130 XA5/XA4/MP3/a_216_n18# XA5/XA4/A 0.15fF
C6131 XA8/XA2/MN1/a_324_n18# XA8/CN1 0.02fF
C6132 XA6/CN0 XA6/CP0 0.59fF
C6133 XA2/CN0 XA2/XA4/A 0.10fF
C6134 XA3/XA12/A XA3/XA9/Y 0.02fF
C6135 XDAC1/XC64a<0>/XRES16/B SARP 21.64fF
C6136 XA3/XA2/MP3/a_216_n18# AVDD 0.07fF
C6137 XA4/XA13/MP1/a_216_n18# XA4/CEO 0.01fF
C6138 XA2/CN1 XA2/XA1/XA1/MN2/S 0.01fF
C6139 XDAC2/XC1/XRES16/B XA0/CN0 0.20fF
C6140 XA2/CN0 XA2/XA5/MN3/a_324_n18# 0.01fF
C6141 XA20/XA3/MN2/a_324_n18# XA20/XA3/N2 0.01fF
C6142 CK_SAMPLE XA20/XA3a/A 0.02fF
C6143 XA2/XA1/XA2/Y XA2/XA1/XA5/MN1/S 0.05fF
C6144 XA3/XA4/MN2/a_324_n18# XA3/XA4/A 0.15fF
C6145 XA1/XA1/XA4/MP1/a_216_n18# XA1/XA1/XA4/MP2/a_216_n18# 0.01fF
C6146 XA3/XA1/XA0/MP1/a_216_n18# XA3/XA1/XA1/MP0/a_216_n18# 0.01fF
C6147 XA3/CN1 AVSS 2.77fF
C6148 XA0/XA5/MP1/a_216_n18# XA0/XA5/MP0/a_216_n18# 0.01fF
C6149 SARN D<8> 0.64fF
C6150 XA1/XA1/XA4/MN2/S AVSS 0.06fF
C6151 XA0/XA4/A XA1/EN 0.11fF
C6152 XA4/XA2/A XA4/XA3/MP0/a_216_n18# 0.08fF
C6153 XB1/XA1/MP0/G AVSS 0.21fF
C6154 XA4/XA2/MP3/a_216_n18# XA4/CN1 0.02fF
C6155 XA20/CPO XA3/XA1/XA1/MP2/a_216_n18# 0.06fF
C6156 XA0/XA3/MP0/a_216_n18# XA0/XA2/MP3/a_216_n18# 0.01fF
C6157 D<1> CK_SAMPLE 0.10fF
C6158 XA3/XA2/MN3/a_324_n18# XA3/CN1 0.03fF
C6159 XA20/XA0/MP1/a_216_n18# AVDD 0.15fF
C6160 XA0/XA9/MP1/a_216_n18# XA0/XA9/MP0/a_216_n18# 0.01fF
C6161 XA6/EN XA5/XA1/XA4/MN0/a_324_n18# 0.07fF
C6162 XB2/XA4/GNG AVDD 4.07fF
C6163 XA4/XA1/XA1/MN2/S XA4/XA1/XA1/MP3/G 0.08fF
C6164 XA5/XA1/XA4/MN1/S XA5/XA1/XA4/MP1/S 0.01fF
C6165 XA8/CEO AVSS 0.26fF
C6166 XA8/CEO XA20/XA12/Y 0.07fF
C6167 XA3/XA11/A XA2/CEO 0.09fF
C6168 XA8/EN XA7/XA9/B 0.07fF
C6169 XA1/XA11/A XA0/CEO 0.09fF
C6170 XA3/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C6171 XA5/CN1 XA5/XA2/MP1/a_216_n18# 0.01fF
C6172 D<2> AVSS 2.25fF
C6173 XA2/XA4/A XA2/XA1/XA4/MN1/S 0.02fF
C6174 XA4/XA2/A D<4> 0.06fF
C6175 XA6/XA9/B XA5/XA9/A 0.02fF
C6176 XA0/CP0 XDAC1/XC0/XRES16/B 0.02fF
C6177 XA0/XA1/XA1/MN0/a_324_n18# XA0/XA1/XA0/MN1/a_324_n18# 0.01fF
C6178 D<1> EN 0.06fF
C6179 XA7/CN0 AVSS 1.26fF
C6180 XA1/XA1/XA1/MN2/S XA20/CNO 0.03fF
C6181 XA4/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C6182 XA1/XA1/XA1/MP3/G XA1/CN1 0.02fF
C6183 XA5/EN XA4/XA4/A 0.11fF
C6184 XA20/XA12/MN0/a_324_n18# DONE 0.06fF
C6185 XDAC2/XC64a<0>/XRES2/B AVSS 3.71fF
C6186 XA0/CP1 XA0/XA3/MN3/a_324_n18# 0.02fF
C6187 XA0/XA5/MP0/a_216_n18# AVDD 0.08fF
C6188 XA2/XA1/XA5/MN2/a_324_n18# XA2/XA2/MN0/a_324_n18# 0.01fF
C6189 XA1/XA13/MN1/a_324_n18# XA1/XA12/MN0/a_324_n18# 0.01fF
C6190 SAR_IN AVDD 0.11fF
C6191 XA1/XA4/A XA1/XA2/A 0.14fF
C6192 VREF XA1/CN0 0.69fF
C6193 XA7/XA11/MP1/a_216_n18# XA7/XA12/MP0/a_216_n18# 0.01fF
C6194 SARP XB1/M4/a_324_n18# 0.01fF
C6195 XA4/XA3/MP2/a_216_n18# XA4/CN1 0.15fF
C6196 XA6/XA9/A XA6/XA9/B 0.29fF
C6197 D<3> AVSS 3.25fF
C6198 XDAC1/XC1/XRES4/B XB1/XA4/GNG 0.16fF
C6199 XA0/CP0 XA0/XA4/MN1/a_324_n18# 0.03fF
C6200 XA8/EN XA7/XA1/XA1/MP3/S 0.10fF
C6201 XA6/XA1/XA5/MN1/a_324_n18# XA20/CNO 0.07fF
C6202 XA3/XA1/XA4/MN2/S XA3/XA1/XA2/Y 0.05fF
C6203 XA6/XA6/MP1/S AVDD 0.12fF
C6204 XA0/XA3/MP3/a_216_n18# XA0/XA3/MP2/a_216_n18# 0.01fF
C6205 XA8/XA2/MN3/a_324_n18# XA8/CN1 0.03fF
C6206 XA8/XA5/MN1/a_324_n18# XA8/CP0 0.15fF
C6207 XA5/XA4/MP3/a_216_n18# VREF 0.03fF
C6208 XA4/XA3/MP3/a_216_n18# VREF 0.03fF
C6209 XA1/XA1/XA5/MN2/a_324_n18# XA1/EN 0.08fF
C6210 XA5/XA9/B XA5/XA9/MN1/a_324_334# 0.07fF
C6211 XA4/XA9/Y XA4/XA11/MP0/a_216_n18# 0.08fF
C6212 XA4/XA1/XA4/MN1/S AVDD 0.02fF
C6213 XA6/XA9/A XA6/XA9/MP1/a_216_n18# 0.08fF
C6214 XDAC2/XC128b<2>/XRES16/B XA0/CN0 0.18fF
C6215 XA7/XA1/XA1/MN2/S AVSS 0.27fF
C6216 XB2/XA0/MP0/a_216_n18# AVDD 0.15fF
C6217 XA6/XA5/MN2/a_324_n18# XA6/XA5/MN1/a_324_n18# 0.01fF
C6218 XB2/XA3/B XDAC2/XC1/XRES2/B 0.05fF
C6219 XA5/XA9/B D<3> 0.05fF
C6220 XA0/XA5/MP2/a_216_n18# XA0/CN0 0.01fF
C6221 XA6/XA1/XA2/MP0/a_216_n18# AVDD 0.08fF
C6222 XA5/XA1/XA4/MN1/a_324_n18# XA5/XA1/XA2/Y 0.09fF
C6223 XA4/XA4/A XA4/XA5/MN0/a_324_n18# 0.07fF
C6224 XA7/XA9/Y XA6/CEO 0.03fF
C6225 XA7/DONE XA7/XA9/B 0.03fF
C6226 XA8/CN1 XA20/XA3a/A 0.01fF
C6227 XDAC2/XC0/XRES1B/B XDAC2/XC0/XRES1A/B 0.01fF
C6228 XDAC1/XC64b<1>/XRES1A/B AVSS 2.95fF
C6229 XDAC2/XC1/XRES2/B AVSS 3.64fF
C6230 XDAC1/XC0/XRES1B/B XDAC1/XC0/XRES16/B 0.13fF
C6231 XDAC2/XC128a<1>/XRES16/B XA0/CN0 0.02fF
C6232 XA0/XA6/MP1/a_216_n18# XA0/XA6/MP0/a_216_n18# 0.01fF
C6233 D<6> XA2/XA2/A 0.06fF
C6234 XA1/XA3/MP2/a_216_n18# XA1/XA3/MP3/a_216_n18# 0.01fF
C6235 XA3/CN0 XA3/XA4/A 0.10fF
C6236 XA7/XA1/XA2/Y XA7/XA2/A 0.01fF
C6237 XA5/XA9/MP1/a_216_334# AVDD 0.09fF
C6238 XA8/CEO CK_SAMPLE 0.09fF
C6239 XA4/XA9/Y XA4/XA9/MN1/a_324_334# 0.09fF
C6240 XA7/XA3/MN3/a_324_n18# XA7/XA4/A 0.01fF
C6241 EN XA3/CN1 0.07fF
C6242 D<2> CK_SAMPLE 0.10fF
C6243 XA4/XA1/XA2/Y XA4/XA1/XA4/MN1/S 0.05fF
C6244 XA8/XA5/MN2/a_324_n18# AVSS 0.01fF
C6245 XA6/XA1/XA5/MN2/S AVDD 0.02fF
C6246 XA3/CP0 XA3/XA4/MN2/a_324_n18# 0.01fF
C6247 XA3/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C6248 XA6/CN0 XA3/CN0 0.30fF
C6249 XA3/XA3/MN3/a_324_n18# XA3/CN1 0.15fF
C6250 XDAC1/XC64b<1>/XRES1A/B XDAC1/X16ab/XRES1B/B 0.63fF
C6251 XDAC2/X16ab/XRES4/B XDAC2/X16ab/XRES8/B 2.60fF
C6252 XA1/XA1/XA4/MP1/S XA1/XA1/XA4/MN1/S 0.01fF
C6253 VREF XA3/EN 1.22fF
C6254 XDAC1/XC32a<0>/XRES1B/B XDAC1/XC128a<1>/XRES16/B 0.05fF
C6255 XA5/XA1/XA5/MN0/a_324_n18# XA5/XA1/XA4/MN2/a_324_n18# 0.01fF
C6256 XA8/XA1/XA1/MP3/G XA20/CPO 0.15fF
C6257 XA7/CN0 CK_SAMPLE 0.08fF
C6258 D<3> XA5/XA3/MN1/a_324_n18# 0.02fF
C6259 XDAC1/X16ab/XRES2/B SARP 3.05fF
C6260 XA2/EN XA2/XA1/XA2/Y 0.14fF
C6261 XA0/XA9/MN1/a_324_n18# XA0/XA9/MN0/a_324_n18# 0.01fF
C6262 XA5/XA1/XA1/MN2/S XA20/CNO 0.03fF
C6263 XA1/XA1/XA4/MP1/a_216_n18# EN 0.15fF
C6264 XA6/XA2/A XA7/XA2/A 0.03fF
C6265 XDAC1/XC64b<1>/XRES8/B SARP 11.94fF
C6266 D<2> EN 0.07fF
C6267 XA3/XA6/MP2/a_216_n18# AVDD 0.09fF
C6268 XA3/XA1/XA1/MP3/S AVDD 0.13fF
C6269 D<3> CK_SAMPLE 0.10fF
C6270 XDAC1/XC128a<1>/XRES16/B XDAC1/XC128a<1>/XRES1B/B 0.12fF
C6271 XA4/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C6272 XA8/EN AVSS 1.45fF
C6273 XA7/CN0 EN 0.06fF
C6274 D<5> XA3/XA6/MP3/a_216_n18# 0.15fF
C6275 XDAC1/XC32a<0>/XRES8/B SARP 11.94fF
C6276 XA2/XA5/MN3/a_324_n18# XA2/XA5/MN2/a_324_n18# 0.01fF
C6277 XA3/XA9/MN1/S AVDD 0.01fF
C6278 XA0/XA5/MP2/a_216_n18# XA0/XA5/MP3/a_216_n18# 0.01fF
C6279 XA6/XA3/MP3/a_216_n18# AVDD 0.07fF
C6280 XA20/XA1/MP0/a_216_334# AVDD 0.16fF
C6281 XB2/XA3/MP0/a_216_334# XB2/XA3/B 0.02fF
C6282 D<3> EN 0.06fF
C6283 XA6/CN0 XA6/XA5/MN1/a_324_n18# 0.02fF
C6284 XA4/XA5/MN1/a_324_n18# XA4/XA5/MN0/a_324_n18# 0.01fF
C6285 XA7/XA13/MN1/a_324_334# AVSS 0.10fF
C6286 XA0/XA1/XA2/Y AVDD 0.33fF
C6287 XDAC1/XC32a<0>/XRES16/B D<4> 0.02fF
C6288 XA5/XA11/MN1/a_324_n18# XA5/XA11/MN0/a_324_n18# 0.01fF
C6289 XA3/XA9/Y XA3/XA9/MN1/S 0.12fF
C6290 XDAC2/XC128b<2>/XRES2/B XDAC2/X16ab/XRES16/B 0.01fF
C6291 XDAC1/XC64a<0>/XRES4/B XDAC1/XC64a<0>/XRES1B/B 1.64fF
C6292 XA6/XA4/A XA6/EN 0.14fF
C6293 XA1/CP0 XA1/XA6/MN0/a_324_n18# 0.07fF
C6294 XB2/XCAPB1/XCAPB3/m3_9828_132# XB2/XA3/B 0.21fF
C6295 XA2/XA6/MP0/a_216_n18# XA2/CN0 0.08fF
C6296 XB1/XA5/MP1/a_216_334# XB1/XA4/GNG 0.01fF
C6297 XA4/XA1/XA5/MN1/S XA4/XA4/A 0.02fF
C6298 XA0/CP1 SARN 0.04fF
C6299 XA4/CEO AVSS 0.49fF
C6300 XA3/XA6/MP0/a_216_n18# AVDD 0.08fF
C6301 XA2/XA8/MP0/a_216_n18# XA2/XA9/A 0.07fF
C6302 XA6/XA4/MP1/a_216_n18# AVDD 0.07fF
C6303 XA1/XA1/XA4/MP1/S XA20/CPO 0.03fF
C6304 XA8/XA1/XA5/MP1/S XA8/XA1/XA5/MP2/S 0.04fF
C6305 XA5/XA11/MN1/a_324_n18# XA5/XA12/MN0/a_324_n18# 0.01fF
C6306 XA1/XA4/A XA1/CN1 0.61fF
C6307 XA20/XA1/MN5/a_324_n18# XA20/XA1/MN6/a_324_n18# 0.01fF
C6308 XA20/CNO XA2/XA1/XA1/MP3/G 0.06fF
C6309 XA7/DONE AVSS 0.15fF
C6310 XA20/XA3/MP1/a_216_n18# AVDD 0.10fF
C6311 D<0> AVSS 0.74fF
C6312 XDAC1/XC1/XRES16/B AVSS 15.88fF
C6313 XA2/XA4/MP0/a_216_n18# XA2/XA4/MP1/a_216_n18# 0.01fF
C6314 XA7/XA4/MP0/a_216_n18# XA7/XA4/MP1/a_216_n18# 0.01fF
C6315 XA6/XA1/XA2/MP0/a_216_n18# XA6/XA1/XA1/MP3/a_216_n18# 0.01fF
C6316 XDAC1/XC0/XRES1A/B SARP 1.50fF
C6317 XA3/CN0 XA3/CP0 4.22fF
C6318 D<5> D<8> 0.04fF
C6319 XA5/XA9/B XA4/CEO 0.02fF
C6320 XA20/XA3/N1 XA20/XA2/MN6/a_324_334# 0.01fF
C6321 XA3/CEO XA2/CEO 0.41fF
C6322 XA4/XA1/XA1/MP3/a_216_n18# XA4/XA1/XA1/MP2/a_216_n18# 0.01fF
C6323 XA5/XA9/MP1/a_216_334# XA5/XA11/MP0/a_216_n18# 0.01fF
C6324 XA0/XA3/MN1/a_324_n18# D<8> 0.16fF
C6325 XA7/XA8/MN0/a_324_n18# XA7/XA7/MN0/a_324_n18# 0.01fF
C6326 XA8/EN CK_SAMPLE 0.09fF
C6327 XA7/XA6/MP3/S XA7/XA9/B 0.07fF
C6328 XA1/XA12/A XA1/XA13/MP1/a_216_n18# 0.08fF
C6329 XA0/CP0 XA1/CN1 0.12fF
C6330 XA7/XA2/MN2/a_324_n18# XA7/CN1 0.02fF
C6331 XA7/XA1/XA1/MN1/a_324_n18# XA20/CNO 0.07fF
C6332 D<5> XA2/XA4/A 0.01fF
C6333 XA2/XA9/Y VREF 0.03fF
C6334 XDAC1/XC1/XRES4/B XDAC1/XC64a<0>/XRES4/B 0.10fF
C6335 XA20/XA1/MN0/a_324_n18# XA20/XA1/MN1/a_324_n18# 0.01fF
C6336 D<4> XA20/CPO 0.06fF
C6337 XB2/XCAPB1/XCAPB0/m3_252_308# XB2/XA4/GNG 0.13fF
C6338 XA8/EN EN 1.01fF
C6339 XA2/XA6/MP0/a_216_n18# XA2/XA5/MP3/a_216_n18# 0.01fF
C6340 XA3/XA5/MN2/a_324_n18# XA3/XA5/MN3/a_324_n18# 0.01fF
C6341 XA5/XA2/MN3/a_324_n18# XA5/XA3/MN0/a_324_n18# 0.01fF
C6342 XA20/XA1/MN4/a_324_n18# XA20/XA1/MP0/S 0.01fF
C6343 XA0/XA3/MP1/a_216_n18# AVDD 0.07fF
C6344 XA8/CN0 XA8/XA6/MP0/a_216_n18# 0.08fF
C6345 XA7/XA9/MP1/a_216_334# XA7/XA9/MP1/a_216_n18# 0.01fF
C6346 XDAC1/XC128b<2>/XRES4/B XDAC1/X16ab/XRES4/B 0.10fF
C6347 XA2/XA1/XA4/MN1/a_324_n18# XA2/XA1/XA4/MN2/a_324_n18# 0.01fF
C6348 XA8/XA12/A DONE 0.02fF
C6349 XDAC1/XC128a<1>/XRES1A/B XDAC1/XC128a<1>/XRES2/B 0.25fF
C6350 XA6/XA6/MN0/a_324_n18# XA6/CP0 0.07fF
C6351 XA8/XA3/MN3/a_324_n18# XA8/CN1 0.15fF
C6352 XA3/XA2/A XA3/EN 0.09fF
C6353 XA0/XA4/A XA0/XA1/XA4/MN2/S 0.06fF
C6354 XDAC1/XC64b<1>/XRES2/B AVSS 3.71fF
C6355 XA8/EN XA8/XA1/XA1/MN2/S 0.05fF
C6356 XA8/XA3/MN2/a_324_n18# AVSS 0.01fF
C6357 XA1/XA13/MP1/a_216_334# XA1/XA13/MP1/a_216_n18# 0.01fF
C6358 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC32a<0>/XRES1B/B 0.03fF
C6359 XA4/XA1/XA5/MP1/S XA20/CNO 0.01fF
C6360 XDAC2/XC32a<0>/XRES8/B AVSS 9.20fF
C6361 XA8/XA1/XA4/MP1/S XA20/CPO 0.03fF
C6362 XA6/XA3/MN0/a_324_n18# XA6/XA3/MN1/a_324_n18# 0.01fF
C6363 XA2/CP0 XA20/CPO 0.05fF
C6364 SAR_IP XB1/XA1/MP0/G 0.01fF
C6365 XDAC1/XC128a<1>/XRES16/B XDAC1/XC128b<2>/XRES16/B 0.41fF
C6366 XA0/XA6/MP1/S VREF 0.04fF
C6367 XA20/CNO XA3/XA4/A 0.21fF
C6368 XA7/XA3/MP3/a_216_n18# VREF 0.03fF
C6369 XA1/XA1/XA1/MP3/G AVSS 0.11fF
C6370 XA4/XA2/MN3/a_324_n18# XA4/CN1 0.03fF
C6371 XB2/M8/a_324_n18# SARN 0.01fF
C6372 XA7/XA1/XA4/MN2/S AVDD 0.02fF
C6373 XA5/CN1 XA5/XA2/A 0.57fF
C6374 XDAC1/XC0/XRES1B/B XA1/CN1 0.01fF
C6375 XDAC1/XC64a<0>/XRES2/B SARP 3.05fF
C6376 XA7/XA1/XA1/MN2/a_324_n18# XA7/XA1/XA1/MN3/a_324_n18# 0.01fF
C6377 XA6/CN0 XA20/CNO 0.06fF
C6378 D<0> CK_SAMPLE 0.11fF
C6379 XA1/XA2/MP1/a_216_n18# XA1/XA2/MP2/a_216_n18# 0.01fF
C6380 XA20/XA12/MP0/a_216_n18# AVDD 0.07fF
C6381 SARN XA20/XA4/MN2/a_324_n18# 0.15fF
C6382 D<1> XA2/CN1 0.04fF
C6383 XA5/XA4/A XA5/XA4/MP0/a_216_n18# 0.07fF
C6384 XA0/XA1/XA1/MN2/S AVDD 0.05fF
C6385 XDAC1/XC128a<1>/XRES4/B XDAC1/XC128b<2>/XRES1A/B 0.01fF
C6386 XA20/XA3/MN2/a_324_n18# XA20/XA3/N1 0.01fF
C6387 XA3/XA1/XA4/MN2/a_324_n18# XA3/XA1/XA5/MN0/a_324_n18# 0.01fF
C6388 XA20/XA3a/MN0/a_324_n18# XA20/XA3/CO 0.07fF
C6389 XA6/CN1 XA6/XA2/MP3/a_216_n18# 0.02fF
C6390 XA6/XA1/XA1/MN2/a_324_n18# XA20/CPO 0.08fF
C6391 XA6/XA1/XA2/Y XA20/CNO 0.22fF
C6392 XA2/XA11/MP1/S XA2/CEO 0.02fF
C6393 XB2/XA0/MP0/a_216_n18# XB2/XA5b/MP1/a_216_n18# 0.01fF
C6394 XA6/XA6/MN2/a_324_n18# AVSS 0.01fF
C6395 XA5/XA2/MP0/a_216_n18# EN 0.08fF
C6396 XA4/XA13/MP1/a_216_n18# XA4/XA12/A 0.08fF
C6397 XA3/XA8/MN0/a_324_n18# XA4/EN 0.06fF
C6398 XA8/XA1/XA5/MP1/S AVDD 0.12fF
C6399 XA0/XA6/MN2/a_324_n18# AVSS 0.01fF
C6400 XA20/XA11/MP1/a_216_n18# XA20/XA11/MP0/a_216_n18# 0.01fF
C6401 XA0/XA5/MP3/a_216_n18# XA0/CN0 0.02fF
C6402 XDAC2/XC64b<1>/XRES16/B SARN 21.64fF
C6403 XA5/CN0 XA5/XA1/XA2/Y 0.02fF
C6404 XA20/XA10/MP1/a_216_n18# AVDD 0.09fF
C6405 XA6/XA5/MP2/a_216_n18# VREF 0.03fF
C6406 XA20/XA9/Y XA20/XA11/Y 0.03fF
C6407 XB2/XA3/MN2/a_324_n18# XB2/XA3/MP0/S 0.09fF
C6408 XA4/CP0 XA4/CN1 0.03fF
C6409 XA8/EN XA7/XA1/XA1/MP2/a_216_n18# 0.02fF
C6410 XDAC1/XC64b<1>/XRES1A/B XDAC1/X16ab/XRES1A/B 0.03fF
C6411 XA20/XA4/MN3/a_324_n18# XA20/XA4/MN2/a_324_n18# 0.01fF
C6412 XA2/EN XA2/XA1/XA5/MN2/a_324_n18# 0.08fF
C6413 XA7/XA3/MN2/a_324_n18# XA7/XA3/MN3/a_324_n18# 0.01fF
C6414 D<0> XA8/XA6/MP3/a_216_n18# 0.15fF
C6415 XA7/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C6416 XA3/XA12/A XA3/XA9/B 0.01fF
C6417 D<2> XA6/XA1/XA1/MP3/G 0.02fF
C6418 XA2/XA9/A XA3/XA9/A 0.01fF
C6419 XA20/XA3/MP3/a_216_n18# XA20/XA3/MP4/a_216_n18# 0.01fF
C6420 XA2/CN0 XA4/EN 0.09fF
C6421 XA7/XA1/XA1/MP3/a_216_n18# XA20/CPO 0.08fF
C6422 XDAC2/XC128b<2>/XRES1A/B AVSS 2.95fF
C6423 XA3/XA1/XA4/MN1/S XA3/XA4/A 0.02fF
C6424 XA0/XA6/MN1/a_324_n18# CK_SAMPLE 0.16fF
C6425 XA20/XA3/MP1/a_216_n18# XA20/XA3/MP2/a_216_n18# 0.01fF
C6426 XA5/XA13/MN1/a_324_334# AVSS 0.10fF
C6427 XA7/XA1/XA1/MN0/a_324_n18# AVSS 0.07fF
C6428 XA6/EN XA4/CP0 0.03fF
C6429 XB1/CKN CK_SAMPLE_BSSW 0.12fF
C6430 XB2/XA4/GNG XDAC2/XC1/XRES1A/B 0.76fF
C6431 XA1/XA1/XA2/MN0/a_324_n18# XA1/XA1/XA4/MN0/a_324_n18# 0.01fF
C6432 XA3/XA1/XA4/MN0/a_324_n18# XA3/XA1/XA2/MN0/a_324_n18# 0.01fF
C6433 XA7/CN1 AVSS 0.80fF
C6434 XA20/XA2/MP6/a_216_334# XA20/XA3/CO 0.15fF
C6435 XA7/XA3/MN2/a_324_n18# XA7/XA4/A 0.01fF
C6436 XA5/XA3/MP0/a_216_n18# XA5/XA2/MP3/a_216_n18# 0.01fF
C6437 XA8/ENO AVSS 0.46fF
C6438 XA0/XA9/MN1/S XA0/XA9/B 0.02fF
C6439 AVDD XA20/XA4/MP6_DMY/a_216_n18# 0.24fF
C6440 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128a<1>/XRES1B/B 0.63fF
C6441 XA6/XA4/A XA6/XA3/MN3/a_324_n18# 0.01fF
C6442 XA3/XA11/A XA3/XA9/A 0.01fF
C6443 XA6/XA4/MP3/a_216_n18# XA6/XA4/A 0.15fF
C6444 XA3/XA1/XA5/MN0/a_324_n18# XA3/XA1/XA2/Y 0.02fF
C6445 XA8/XA5/MP2/a_216_n18# XA8/XA5/MP1/a_216_n18# 0.01fF
C6446 XA0/CP1 XA0/XA6/MP1/a_216_n18# 0.01fF
C6447 XA4/XA1/XA4/MN2/S AVDD 0.02fF
C6448 XA3/XA1/XA4/MN2/S XA3/XA1/XA4/MP2/S 0.01fF
C6449 XA1/XA4/A XA1/XA4/MN2/a_324_n18# 0.15fF
C6450 XA2/CN1 XA3/CN1 2.07fF
C6451 XDAC1/XC64b<1>/XRES2/B XDAC1/XC0/XRES2/B 0.05fF
C6452 XA0/XA6/MP0/a_216_n18# AVDD 0.08fF
C6453 XA20/XA9/A XA20/XA11/Y 0.25fF
C6454 XA1/XA1/XA2/Y AVDD 0.33fF
C6455 XA1/XA1/XA5/MP1/S AVDD 0.13fF
C6456 XA6/XA1/XA4/MP1/S EN 0.02fF
C6457 D<6> XA0/CN0 0.05fF
C6458 XA0/XA4/A XA0/CN0 0.10fF
C6459 XA5/XA2/A XA5/XA2/MN0/a_324_n18# 0.08fF
C6460 D<0> XA8/CN1 0.38fF
C6461 XA1/XA1/XA1/MP3/G EN 0.10fF
C6462 XA3/XA6/MP3/a_216_n18# AVDD 0.08fF
C6463 XA5/XA4/MP0/a_216_n18# VREF 0.02fF
C6464 XA3/CP0 XA20/CNO 0.05fF
C6465 D<2> XA2/CN1 0.04fF
C6466 XA1/XA9/Y XA0/CEO 0.03fF
C6467 XDAC2/XC1/XRES1A/B XDAC2/XC64a<0>/XRES1A/B 0.03fF
C6468 D<5> XA0/CP1 0.22fF
C6469 XA4/XA1/XA2/Y XA4/XA1/XA4/MN2/S 0.05fF
C6470 XA6/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C6471 XA7/XA11/MP0/a_216_n18# XA7/XA9/Y 0.08fF
C6472 XA20/XA3a/A XA20/XA2a/MP2/a_216_n18# 0.01fF
C6473 XA4/XA2/MN1/a_324_n18# XA4/CN1 0.02fF
C6474 XA1/CP0 D<4> 0.11fF
C6475 XA6/XA1/XA5/MN1/S AVSS 0.12fF
C6476 XA6/XA9/B XA6/DONE 0.03fF
C6477 XA0/XA6/MN2/a_324_n18# CK_SAMPLE 0.15fF
C6478 XA4/XA1/XA1/MP3/G XA4/XA1/XA2/MN0/a_324_n18# 0.06fF
C6479 XA7/CN0 XA2/CN1 0.09fF
C6480 XA2/CN0 SARN 0.08fF
C6481 XA2/XA9/MN1/a_324_334# XA2/XA11/MN0/a_324_n18# 0.01fF
C6482 XA0/CP1 XA0/XA3/MN1/a_324_n18# 0.02fF
C6483 XA4/XA3/MN1/a_324_n18# XA4/XA3/MN2/a_324_n18# 0.01fF
C6484 XA1/XA6/MN3/S AVDD 0.01fF
C6485 XB2/XCAPB1/XCAPB0/m3_9828_132# XB2/XA3/B 0.21fF
C6486 XA8/CN0 AVSS 0.56fF
C6487 XA2/XA11/MP0/a_216_n18# XA2/XA11/MP1/a_216_n18# 0.01fF
C6488 XA2/XA1/XA1/MP0/a_216_n18# XA3/EN 0.01fF
C6489 XA1/XA3/MN3/a_324_n18# XA1/CN1 0.15fF
C6490 CK_SAMPLE_BSSW XB1/XA3/MN0/a_324_n18# 0.07fF
C6491 XA8/XA1/XA5/MN1/S AVDD 0.02fF
C6492 XA8/XA3/MP3/a_216_n18# XA8/XA4/MP0/a_216_n18# 0.01fF
C6493 D<3> XA2/CN1 0.03fF
C6494 XA0/XA1/XA1/MP3/G AVDD 0.63fF
C6495 XDAC2/XC128b<2>/XRES16/B XDAC2/X16ab/XRES16/B 0.41fF
C6496 XA7/XA2/MP0/a_216_n18# EN 0.08fF
C6497 XA7/XA4/A XA7/EN 0.20fF
C6498 XA8/XA4/MP0/a_216_n18# XA8/XA4/MP1/a_216_n18# 0.01fF
C6499 XA2/XA9/B XA2/XA9/MP1/a_216_334# 0.08fF
C6500 XA6/XA5/MN0/a_324_n18# XA6/CP0 0.09fF
C6501 XA7/CEO XA8/XA11/A 0.08fF
C6502 XA5/XA5/MP1/a_216_n18# AVDD 0.07fF
C6503 D<6> XA2/XA3/MP3/a_216_n18# 0.02fF
C6504 XA2/XA5/MP3/a_216_n18# XA2/CN0 0.02fF
C6505 XA5/XA13/MN1/a_324_n18# XA5/XA12/MN0/a_324_n18# 0.01fF
C6506 XA8/ENO CK_SAMPLE 0.13fF
C6507 XA7/XA1/XA4/MN1/a_324_n18# XA7/XA1/XA4/MN2/a_324_n18# 0.01fF
C6508 XDAC2/XC128a<1>/XRES4/B AVSS 5.49fF
C6509 XA0/CN0 SARP 0.02fF
C6510 XA2/CP0 XA1/CP0 1.65fF
C6511 XDAC1/X16ab/XRES4/B AVSS 5.49fF
C6512 XA8/XA1/XA4/MP2/S AVDD 0.11fF
C6513 XB1/XA2/MP0/G XB1/XA4/GNG 0.07fF
C6514 XA8/XA3/MN2/a_324_n18# XA8/CN1 0.16fF
C6515 XA8/XA3/MP2/a_216_n18# AVDD 0.07fF
C6516 XA7/XA1/XA2/Y XA7/XA1/XA5/MN1/a_324_n18# 0.08fF
C6517 XA7/XA2/MP3/a_216_n18# XA7/CN1 0.02fF
C6518 XA8/XA6/MN2/a_324_n18# XA8/XA6/MN1/a_324_n18# 0.01fF
C6519 XDAC2/X16ab/XRES1A/B XDAC2/X16ab/XRES1B/B 0.01fF
C6520 XA8/XA1/XA1/MP1/a_216_n18# XA20/CNO 0.06fF
C6521 XA20/XA9/MN0/a_324_334# XA20/XA9/MN0/a_324_n18# 0.01fF
C6522 VREF XA20/XA3a/A 0.20fF
C6523 XDAC1/XC1/XRES1A/B AVSS 2.78fF
C6524 XA1/XA4/A AVSS 1.07fF
C6525 XA5/XA7/MN0/a_324_n18# XA5/XA6/MN3/a_324_n18# 0.01fF
C6526 XA6/XA4/MN0/a_324_n18# AVSS 0.01fF
C6527 XA8/EN XA6/XA1/XA1/MP3/G 0.01fF
C6528 XA5/XA2/MN0/a_324_n18# XA5/XA1/XA5/MN2/a_324_n18# 0.01fF
C6529 XA4/XA4/MP0/a_216_n18# XA4/XA4/A 0.07fF
C6530 D<7> XA3/CN1 0.13fF
C6531 XA7/CN1 EN 0.02fF
C6532 AVDD D<8> 1.41fF
C6533 XA3/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C6534 XDAC2/XC128a<1>/XRES1B/B XDAC2/XC128a<1>/XRES4/B 1.64fF
C6535 XDAC2/XC128a<1>/XRES2/B XDAC2/XC128a<1>/XRES8/B 1.58fF
C6536 XA8/ENO EN 0.74fF
C6537 XA2/XA5/MP1/a_216_n18# AVDD 0.07fF
C6538 XDAC2/XC1/XRES16/B XDAC2/XC1/XRES8/B 1.42fF
C6539 XDAC1/X16ab/XRES1B/B XDAC1/X16ab/XRES4/B 1.64fF
C6540 XDAC1/X16ab/XRES2/B XDAC1/X16ab/XRES8/B 1.58fF
C6541 XA3/CEO XA4/XA11/MP1/a_216_n18# 0.06fF
C6542 XA5/XA1/XA1/MP3/G D<3> 0.02fF
C6543 XA1/CP0 XA1/XA4/MP1/a_216_n18# 0.02fF
C6544 D<1> VREF 1.75fF
C6545 XA0/XA9/B XA1/EN 0.07fF
C6546 XDAC2/XC1/XRES1B/B SARN 1.79fF
C6547 XA0/XA2/MP1/a_216_n18# D<8> 0.02fF
C6548 XDAC1/XC64b<1>/XRES8/B XDAC1/X16ab/XRES8/B 0.21fF
C6549 XA0/CP0 AVSS 2.25fF
C6550 XA4/XA1/XA2/Y XA4/XA1/XA4/MN2/a_324_n18# 0.08fF
C6551 XA5/XA6/MN3/S AVSS 0.13fF
C6552 XA6/XA9/MP1/a_216_n18# XA6/XA9/MP0/a_216_n18# 0.01fF
C6553 SARN XA20/XA4/MN3/a_324_n18# 0.15fF
C6554 XA2/XA4/A AVDD 1.42fF
C6555 XA5/XA9/A XA5/XA8/MN0/a_324_n18# 0.09fF
C6556 XA4/XA4/MP3/a_216_n18# XA4/XA5/MP0/a_216_n18# 0.01fF
C6557 XDAC1/XC64b<1>/XRES4/B XDAC1/XC64b<1>/XRES16/B 0.25fF
C6558 XA20/CPO XA1/CN0 0.06fF
C6559 XA8/ENO XA8/XA1/XA1/MN2/S 0.06fF
C6560 XA6/XA6/MN1/S AVSS 0.15fF
C6561 XA20/XA3a/MP1/a_216_n18# XA20/XA3a/MP2/a_216_n18# 0.01fF
C6562 XB2/XA3/B XB2/XA4/MP1/a_216_n18# 0.01fF
C6563 XA4/XA1/XA1/MP3/G XA20/CPO 0.14fF
C6564 XA2/XA1/XA4/MP0/a_216_n18# XA2/XA1/XA4/MP1/a_216_n18# 0.01fF
C6565 XA5/XA2/A XA5/XA2/MN1/a_324_n18# 0.15fF
C6566 XA0/XA4/MP2/a_216_n18# XA0/XA4/MP1/a_216_n18# 0.01fF
C6567 XA6/XA6/MP3/S XA7/EN 0.02fF
C6568 XA6/XA4/MN3/a_324_n18# XA6/XA4/MN2/a_324_n18# 0.01fF
C6569 CK_SAMPLE XA8/CN0 0.04fF
C6570 XA4/XA11/MP1/S AVDD 0.19fF
C6571 XA7/CP0 AVDD 1.31fF
C6572 XA5/XA1/XA4/MP2/a_216_n18# XA5/XA1/XA4/MP1/a_216_n18# 0.01fF
C6573 XDAC2/XC64a<0>/XRES1B/B XDAC2/XC64a<0>/XRES4/B 1.64fF
C6574 XA5/XA9/B XA5/XA6/MN3/S 0.09fF
C6575 XA1/XA12/MP0/a_216_n18# AVDD 0.08fF
C6576 XA6/XA1/XA4/MN0/a_324_n18# XA7/EN 0.07fF
C6577 D<3> XA5/XA4/A 0.26fF
C6578 XA1/XA1/XA2/MN0/a_324_n18# XA1/XA1/XA1/MN3/a_324_n18# 0.01fF
C6579 XA6/XA1/XA5/MN1/S EN 0.01fF
C6580 XDAC1/XC1/XRES1B/B SARP 1.79fF
C6581 XA5/XA9/B XA5/XA6/MP1/S 0.07fF
C6582 D<7> D<3> 0.01fF
C6583 XA6/XA9/B XA6/XA11/A 0.03fF
C6584 XA6/XA4/MP0/a_216_n18# XA6/XA3/MP3/a_216_n18# 0.01fF
C6585 XDAC1/XC32a<0>/XRES4/B XDAC1/XC32a<0>/XRES16/B 0.25fF
C6586 XA7/XA12/A XA7/XA13/MN1/a_324_n18# 0.07fF
C6587 XA4/XA12/A AVSS 0.42fF
C6588 XA6/XA1/XA5/MP2/S XA6/XA1/XA5/MP1/S 0.04fF
C6589 XA6/XA1/XA1/MP0/a_216_n18# XA6/XA1/XA0/MP1/a_216_n18# 0.01fF
C6590 XA3/XA11/MP1/a_216_n18# XA2/CEO 0.07fF
C6591 XA3/XA3/MP1/a_216_n18# XA3/CN1 0.15fF
C6592 EN XA2/XA1/XA4/MP1/S 0.02fF
C6593 XA3/XA9/B XA3/XA9/MN1/S 0.02fF
C6594 XA7/XA6/MP0/a_216_n18# XA7/XA6/MP1/a_216_n18# 0.01fF
C6595 XA0/XA9/B XA0/DONE 0.03fF
C6596 XA4/CN1 AVDD 1.31fF
C6597 XA7/CN1 XA8/CN1 0.10fF
C6598 XA8/XA11/A XA8/XA11/MN0/a_324_n18# 0.09fF
C6599 AVDD XA7/XA3/MP0/a_216_n18# 0.08fF
C6600 XA1/XA2/A XA1/XA3/MN0/a_324_n18# 0.07fF
C6601 XA8/EN XA8/XA1/XA1/MN0/a_324_n18# 0.08fF
C6602 XA5/XA9/Y XA5/XA11/A 0.14fF
C6603 XA8/ENO XA8/CN1 0.10fF
C6604 XDAC1/XC0/XRES1B/B AVSS 2.91fF
C6605 AVDD XA2/XA1/XA4/MP1/a_216_n18# 0.08fF
C6606 VREF XA3/CN1 0.77fF
C6607 XB2/XA5/MP1/a_216_n18# AVDD 0.13fF
C6608 VREF XA1/XA5/MP2/a_216_n18# 0.03fF
C6609 XA20/CPO XA3/EN 0.63fF
C6610 XDAC1/XC128a<1>/XRES2/B XDAC1/XC128b<2>/XRES2/B 0.05fF
C6611 XA3/DONE AVDD 0.21fF
C6612 XA4/XA2/A XA4/XA1/XA5/MN2/S 0.05fF
C6613 XA6/EN AVDD 4.07fF
C6614 XA8/XA4/MN2/a_324_n18# AVSS 0.01fF
C6615 XA6/XA4/MP0/a_216_n18# XA6/XA4/MP1/a_216_n18# 0.01fF
C6616 XA0/CP1 XA0/XA9/A 0.01fF
C6617 XA0/XA2/MP0/a_216_n18# AVDD 0.08fF
C6618 XA2/XA7/MN0/a_324_n18# XA2/XA8/MN0/a_324_n18# 0.01fF
C6619 XA7/XA1/XA2/Y AVSS 0.31fF
C6620 XA5/XA9/MP1/a_216_n18# XA5/XA9/MP1/a_216_334# 0.01fF
C6621 XA20/CNO XA20/XA3/CO 0.76fF
C6622 XA8/CEO VREF 0.18fF
C6623 XA1/XA4/A EN 0.09fF
C6624 XA0/CP0 CK_SAMPLE 0.09fF
C6625 XA5/XA1/XA5/MN1/S XA20/CNO 0.01fF
C6626 XA7/XA13/MP1/a_216_n18# XA7/XA13/MP1/a_216_334# 0.01fF
C6627 XA5/XA6/MN3/S CK_SAMPLE 0.03fF
C6628 XDAC2/XC128a<1>/XRES1A/B XDAC2/XC32a<0>/XRES1B/B 0.63fF
C6629 XB2/XA5/MN1/a_324_334# XB2/XA5/MN1/a_324_n18# 0.01fF
C6630 XA5/XA12/A AVDD 0.44fF
C6631 D<2> VREF 1.75fF
C6632 XDAC1/XC64b<1>/XRES4/B XDAC1/XC0/XRES8/B 0.01fF
C6633 XA4/XA12/MN0/a_324_n18# AVSS 0.01fF
C6634 XDAC1/XC32a<0>/XRES4/B XDAC1/XC32a<0>/XRES2/B 0.55fF
C6635 XA0/XA2/MP0/a_216_n18# XA0/XA2/MP1/a_216_n18# 0.01fF
C6636 XA2/EN XA2/XA1/XA4/MN2/S 0.02fF
C6637 XA4/XA4/A AVSS 1.10fF
C6638 XA5/XA6/MP1/S CK_SAMPLE 0.02fF
C6639 XA3/XA9/Y XA3/DONE 0.06fF
C6640 XA6/XA6/MN1/S CK_SAMPLE 0.04fF
C6641 XA3/XA1/XA4/MN1/a_324_n18# XA20/CPO 0.08fF
C6642 XDAC1/XC128a<1>/XRES8/B XDAC1/XC128a<1>/XRES16/B 1.42fF
C6643 XA4/XA6/MP3/S AVDD 0.16fF
C6644 XA1/XA1/XA5/MN1/S AVSS 0.12fF
C6645 XA7/CN0 VREF 0.69fF
C6646 D<6> SARP 0.12fF
C6647 XA6/XA11/MP1/a_216_n18# AVDD 0.08fF
C6648 XA2/EN XA1/XA1/XA1/MP2/S 0.14fF
C6649 XA3/XA1/XA4/MN0/a_324_n18# XA20/CPO 0.09fF
C6650 XA3/XA6/MP1/a_216_n18# XA3/XA6/MP2/a_216_n18# 0.01fF
C6651 XA0/CP0 EN 0.08fF
C6652 XA20/XA9/Y SARN 0.66fF
C6653 XA6/XA2/A AVSS 0.28fF
C6654 XA3/XA9/MP1/a_216_334# AVDD 0.09fF
C6655 XA6/XA3/MN0/a_324_n18# XA6/CN1 0.10fF
C6656 XA5/CEO XA6/XA12/MN0/a_324_n18# 0.07fF
C6657 XA4/XA11/A AVSS 0.28fF
C6658 XA3/XA1/XA5/MP1/a_216_n18# AVDD 0.08fF
C6659 XA4/XA1/XA5/MN1/a_324_n18# XA4/XA1/XA5/MN0/a_324_n18# 0.01fF
C6660 D<5> XA4/EN 0.45fF
C6661 XB2/XCAPB1/XCAPB1/m3_9756_132# XB2/XA4/GNG 0.02fF
C6662 XA0/XA1/XA1/MN1/a_324_n18# XA0/XA1/XA1/MN2/a_324_n18# 0.01fF
C6663 XB2/XA3/B CK_SAMPLE_BSSW 0.05fF
C6664 XA20/XA2/MP3/a_216_n18# XA20/XA9/Y 0.07fF
C6665 D<3> VREF 1.75fF
C6666 XA20/XA3/N2 XA20/XA3a/A 0.07fF
C6667 XB1/XA4/MN1/S AVSS 0.14fF
C6668 XA5/XA2/A XA5/CN0 0.05fF
C6669 XA6/XA5/MP1/a_216_n18# XA6/CP0 0.15fF
C6670 XA6/XA1/XA4/MP2/S XA6/XA4/A 0.05fF
C6671 XA5/XA5/MP2/a_216_n18# XA5/XA5/MP3/a_216_n18# 0.01fF
C6672 XA2/XA11/MN0/a_324_n18# XA2/XA11/A 0.09fF
C6673 XA3/XA9/MP1/a_216_334# XA3/XA9/Y 0.07fF
C6674 XA4/XA1/XA1/MP3/G XA4/XA1/XA1/MP1/a_216_n18# 0.01fF
C6675 XA0/XA4/A XA0/XA5/MN0/a_324_n18# 0.07fF
C6676 CK_SAMPLE_BSSW AVSS 0.83fF
C6677 XA8/XA4/MP3/a_216_n18# AVDD 0.07fF
C6678 XDAC2/XC128b<2>/XRES16/B XDAC2/XC128a<1>/XRES8/B 0.03fF
C6679 XA3/XA1/XA4/MP1/S XA4/EN 0.02fF
C6680 XDAC2/X16ab/XRES16/B XA0/CN0 0.03fF
C6681 XA0/XA1/XA5/MN2/S AVDD 0.02fF
C6682 XA20/XA1/MP4_DMY/a_216_n18# XA20/XA1/MP5_DMY/a_216_n18# 0.01fF
C6683 XA8/XA1/XA4/MN1/a_324_n18# XA8/XA1/XA2/Y 0.09fF
C6684 XA20/XA3a/A XA8/CP0 0.01fF
C6685 XA2/XA6/MP1/S D<6> 0.02fF
C6686 XA3/XA3/MN1/a_324_n18# XA3/XA3/MN0/a_324_n18# 0.01fF
C6687 XDAC2/XC128b<2>/XRES1B/B SARN 1.79fF
C6688 XA2/CN1 XA2/XA2/MN3/a_324_n18# 0.03fF
C6689 XA6/XA5/MN0/a_324_n18# XA6/XA5/MN1/a_324_n18# 0.01fF
C6690 XA5/CN1 XA5/XA2/MN1/a_324_n18# 0.02fF
C6691 XA20/XA3a/A XA20/XA4/MN0/a_324_n18# 0.06fF
C6692 XA5/XA1/XA5/MP2/a_216_n18# AVDD 0.08fF
C6693 XA8/XA1/XA1/MP0/a_216_n18# EN 0.06fF
C6694 XA4/EN XA3/XA1/XA1/MN2/S 0.12fF
C6695 EN XA0/XA1/XA1/MN1/a_324_n18# 0.07fF
C6696 XB2/M6/a_324_n18# XB2/M5/a_324_n18# 0.01fF
C6697 XA7/XA1/XA5/MN1/a_324_n18# XA7/XA1/XA5/MN2/a_324_n18# 0.01fF
C6698 D<5> XA2/CN0 0.06fF
C6699 XA7/XA1/XA4/MN1/a_324_n18# XA7/XA1/XA4/MN0/a_324_n18# 0.01fF
C6700 XA3/XA3/MN2/a_324_n18# XA3/XA4/A 0.01fF
C6701 XDAC1/XC64a<0>/XRES16/B XDAC1/XC64a<0>/XRES4/B 0.25fF
C6702 XA4/CN0 XA0/CN0 0.13fF
C6703 XDAC2/XC128a<1>/XRES8/B XDAC2/XC128a<1>/XRES16/B 1.42fF
C6704 XA8/XA11/A AVSS 0.28fF
C6705 XA6/XA6/MP1/a_216_n18# XA6/XA6/MP0/a_216_n18# 0.01fF
C6706 XA20/XA9/A SARN 1.02fF
C6707 XA5/XA2/MP3/a_216_n18# VREF 0.03fF
C6708 XA3/XA1/XA1/MP3/S XA3/XA1/XA1/MP3/G 0.04fF
C6709 XA7/XA1/XA0/MN1/a_324_n18# AVSS 0.09fF
C6710 XA3/XA12/A AVSS 0.39fF
C6711 XA7/XA5/MN0/a_324_n18# XA7/XA4/MN3/a_324_n18# 0.01fF
C6712 XA5/XA9/Y XA5/CEO 0.03fF
C6713 XA3/XA6/MP0/a_216_n18# XA3/XA6/MP1/a_216_n18# 0.01fF
C6714 XA5/CN0 XA0/CN0 0.13fF
C6715 XA1/XA1/XA2/Y XA1/XA2/A 0.01fF
C6716 XA4/XA4/MP3/a_216_n18# VREF 0.03fF
C6717 VREF XA8/XA6/MP1/a_216_n18# 0.01fF
C6718 XA4/XA5/MP2/a_216_n18# XA4/CP0 0.15fF
C6719 XA0/CP1 AVDD 1.85fF
C6720 XDAC1/XC0/XRES1A/B XDAC1/XC0/XRES4/B 0.29fF
C6721 XDAC1/XC0/XRES2/B XDAC1/XC0/XRES1B/B 0.23fF
C6722 XB1/XCAPB1/XCAPB1/m3_9756_132# XB1/XA3/B 0.07fF
C6723 XB1/XA3/MP2/a_216_n18# XB1/XA4/GNG 0.02fF
C6724 XA20/XA11/Y AVDD 0.48fF
C6725 XA1/CP0 XA1/CN0 4.42fF
C6726 XB1/XA5/MP1/a_216_n18# XB1/XA5/MP1/a_216_334# 0.01fF
C6727 XA5/XA5/MP3/a_216_n18# VREF 0.02fF
C6728 XA1/XA8/MN0/a_324_n18# XA1/XA9/A 0.09fF
C6729 D<5> SARN 0.03fF
C6730 XA0/CP0 XA0/XA4/MN2/a_324_n18# 0.01fF
C6731 XA4/XA1/XA1/MP0/a_216_n18# XA4/XA1/XA1/MP1/a_216_n18# 0.01fF
C6732 XA20/CNO XA1/EN 0.93fF
C6733 XA7/XA1/XA2/Y EN 0.07fF
C6734 XA2/XA1/XA5/MP2/a_216_n18# XA2/XA2/MP0/a_216_n18# 0.01fF
C6735 XDAC2/XC1/XRES16/B XDAC2/XC64a<0>/XRES16/B 0.41fF
C6736 XA5/CEO XA5/XA11/A 0.05fF
C6737 D<0> XA8/XA9/B 0.05fF
C6738 XA0/CP1 XDAC1/XC128b<2>/XRES16/B 0.05fF
C6739 XA0/XA6/MN1/a_324_n18# XA0/XA6/MN0/a_324_n18# 0.01fF
C6740 XA3/XA5/MN2/a_324_n18# AVSS 0.01fF
C6741 XA4/XA4/A EN 0.10fF
C6742 XA3/XA5/MP2/a_216_n18# XA3/XA5/MP1/a_216_n18# 0.01fF
C6743 XA7/XA1/XA4/MP2/a_216_n18# XA7/XA1/XA5/MP0/a_216_n18# 0.01fF
C6744 XB2/XA4/GNG XB2/XA3/B 434.15fF
C6745 XA5/XA1/XA4/MP2/a_216_n18# EN 0.15fF
C6746 XA5/EN XA4/CN1 0.10fF
C6747 XDAC2/XC0/XRES2/B SARN 3.08fF
C6748 XA2/XA6/MP0/a_216_n18# AVDD 0.08fF
C6749 XA6/XA1/XA5/MP0/a_216_n18# XA6/XA1/XA4/MP2/a_216_n18# 0.01fF
C6750 XA2/EN XA1/XA9/B 0.07fF
C6751 XA5/XA3/MN2/a_324_n18# AVSS 0.01fF
C6752 XA1/XA1/XA5/MN1/S EN 0.01fF
C6753 XA2/XA12/A XA2/XA12/MP0/a_216_n18# 0.07fF
C6754 XA8/EN VREF 1.22fF
C6755 XA8/XA2/MP2/a_216_n18# XA8/XA2/A 0.15fF
C6756 XA2/XA11/MN0/a_324_n18# AVSS 0.01fF
C6757 XA6/XA1/XA4/MP2/a_216_n18# AVDD 0.08fF
C6758 XA0/XA12/A XA0/XA11/MP1/S 0.06fF
C6759 XB2/XA4/GNG AVSS 5.22fF
C6760 XA7/XA2/MP2/a_216_n18# AVDD 0.07fF
C6761 XDAC1/X16ab/XRES1A/B XDAC1/X16ab/XRES4/B 0.29fF
C6762 XA1/XA1/XA5/MP2/S AVDD 0.08fF
C6763 XA6/XA2/A EN 0.13fF
C6764 XA20/XA11/MP1/S DONE 0.02fF
C6765 D<0> XA8/XA6/MP3/S 0.02fF
C6766 XA3/XA2/A XA3/CN1 0.63fF
C6767 XA1/XA3/MN0/a_324_n18# XA1/CN1 0.10fF
C6768 XA6/EN XA5/EN 1.82fF
C6769 XA2/XA4/MN3/a_324_n18# XA2/XA5/MN0/a_324_n18# 0.01fF
C6770 XA1/XA6/MP2/a_216_n18# XA1/XA6/MP3/a_216_n18# 0.01fF
C6771 XA3/XA12/MN0/a_324_n18# XA2/CEO 0.07fF
C6772 XA8/XA1/XA1/MP2/a_216_n18# AVDD 0.08fF
C6773 XA1/XA1/XA5/MP2/S XA1/XA1/XA5/MN2/S 0.01fF
C6774 XDAC2/X16ab/XRES2/B XDAC2/X16ab/XRES16/B 1.61fF
C6775 SAR_IN XB2/XA3/B 0.23fF
C6776 XA3/EN XA2/XA1/XA1/MP3/S 0.10fF
C6777 XA4/DONE XA4/XA9/B 0.03fF
C6778 XA4/XA6/MP3/S XA5/EN 0.02fF
C6779 XA8/EN XA7/XA1/XA1/MP2/S 0.14fF
C6780 XA3/XA4/MP0/a_216_n18# XA3/CN1 0.08fF
C6781 XA5/XA2/MN1/a_324_n18# XA5/XA2/MN0/a_324_n18# 0.01fF
C6782 XB2/XA0/MN0/a_324_n18# CK_SAMPLE_BSSW 0.08fF
C6783 XA1/XA1/XA5/MP2/a_216_n18# EN 0.16fF
C6784 XA5/CN1 XA5/CN0 0.09fF
C6785 XA6/EN XA5/XA1/XA2/MP0/a_216_n18# 0.08fF
C6786 XDAC2/XC64b<1>/XRES1A/B XDAC2/X16ab/XRES4/B 0.01fF
C6787 XA3/CN0 XA3/XA1/XA2/Y 0.02fF
C6788 SAR_IN AVSS 0.78fF
C6789 XA7/XA5/MP3/a_216_n18# XA7/XA5/MP2/a_216_n18# 0.01fF
C6790 SAR_IN XB2/M5/a_324_n18# 0.02fF
C6791 XDAC2/XC1/XRES4/B XDAC2/XC1/XRES1A/B 0.29fF
C6792 XA0/XA1/XA5/MP2/a_216_n18# XA0/XA2/MP0/a_216_n18# 0.01fF
C6793 XA1/XA11/A XA1/XA12/A 0.07fF
C6794 XA7/XA4/MP0/a_216_n18# XA7/XA4/A 0.07fF
C6795 XA6/XA4/MN1/a_324_n18# XA6/XA4/A 0.15fF
C6796 XA1/XA9/B XA1/XA9/MN0/a_324_n18# 0.01fF
C6797 XA5/XA1/XA2/Y XA20/CNO 0.22fF
C6798 XA2/XA1/XA5/MN2/S AVDD 0.02fF
C6799 XA3/XA3/MN0/a_324_n18# XA3/CN1 0.10fF
C6800 XA4/CEO VREF 0.23fF
C6801 XA20/XA2/MN1/a_324_n18# SARP 0.09fF
C6802 XA0/XA11/A XA0/XA11/MP1/a_216_n18# 0.08fF
C6803 XDAC2/XC1/XRES8/B XA0/CN0 0.01fF
C6804 XA0/XA1/XA4/MN1/S AVDD 0.02fF
C6805 XA6/XA1/XA1/MN1/a_324_n18# XA6/XA1/XA1/MN0/a_324_n18# 0.01fF
C6806 XDAC2/XC64a<0>/XRES1A/B AVSS 2.97fF
C6807 XB2/XA0/MP0/a_216_n18# XB2/XA3/B 0.01fF
C6808 AVDD XA2/XA2/MP0/a_216_n18# 0.08fF
C6809 XA6/XA4/MP3/a_216_n18# AVDD 0.07fF
C6810 XA5/XA3/MP2/a_216_n18# VREF 0.03fF
C6811 XB2/XA4/MP0/a_216_n18# AVDD 0.09fF
C6812 XA5/XA3/MN2/a_324_n18# XA5/XA3/MN1/a_324_n18# 0.01fF
C6813 D<7> XA1/XA1/XA1/MP3/G 0.02fF
C6814 XA8/EN XA8/XA1/XA2/Y 0.14fF
C6815 XA4/XA1/XA4/MN1/S AVSS 0.10fF
C6816 XA2/XA4/A XA1/XA2/A 0.03fF
C6817 XB1/XCAPB1/XCAPB0/m3_9828_132# XB1/XA4/GNG 0.03fF
C6818 XA7/XA3/MP0/a_216_n18# XA7/XA2/A 0.08fF
C6819 XA7/XA1/XA1/MP3/G XA7/XA1/XA1/MP3/a_216_n18# 0.07fF
C6820 XB2/M4/a_324_n18# SARN 0.01fF
C6821 D<0> VREF 1.60fF
C6822 XA3/XA2/MP2/a_216_n18# AVDD 0.07fF
C6823 XA2/EN XA1/XA1/XA4/MP1/S 0.02fF
C6824 XA2/XA2/A XA20/CNO 0.03fF
C6825 XA3/XA1/XA5/MN1/S XA20/CNO 0.01fF
C6826 XA20/XA0/MN1/a_324_n18# AVSS 0.09fF
C6827 XB1/XA3/MP0/a_216_n18# XB1/XA4/GNG 0.01fF
C6828 XA4/XA9/A XA4/XA11/A 0.01fF
C6829 XA0/CEIN XB1/XA3/B 0.02fF
C6830 XA3/XA1/XA5/MP1/S XA20/CNO 0.01fF
C6831 XDAC2/XC64b<1>/XRES2/B XDAC2/XC64b<1>/XRES16/B 1.61fF
C6832 XA20/XA9/Y XA20/XA9/A 2.03fF
C6833 XA4/XA2/A XA3/CN1 0.04fF
C6834 XA0/CEIN XB1/M5/a_324_n18# 0.08fF
C6835 XDAC2/XC64a<0>/XRES8/B XDAC2/XC64a<0>/XRES2/B 1.58fF
C6836 XB1/M7/a_324_n18# SARP 0.02fF
C6837 XA4/XA5/MN2/a_324_n18# AVSS 0.01fF
C6838 XB2/CKN XB2/XA3/MN1/a_324_n18# 0.15fF
C6839 XA6/XA1/XA5/MN2/S AVSS 0.09fF
C6840 XA4/XA5/MP2/a_216_n18# XA4/XA5/MP1/a_216_n18# 0.01fF
C6841 XA4/XA9/Y XA3/CEO 0.01fF
C6842 XDAC1/XC32a<0>/XRES8/B XDAC1/XC64a<0>/XRES4/B 0.01fF
C6843 XDAC2/XC128b<2>/XRES1A/B XDAC2/XC128b<2>/XRES8/B 0.12fF
C6844 XDAC2/XC128b<2>/XRES2/B XDAC2/XC128b<2>/XRES4/B 0.55fF
C6845 XA20/XA2/MP0/a_216_n18# XA20/XA1/MP6_DMY/a_216_n18# 0.01fF
C6846 XA6/XA6/MP1/a_216_n18# AVDD 0.08fF
C6847 XA8/XA1/XA1/MP2/a_216_n18# XA8/XA1/XA1/MP3/a_216_n18# 0.01fF
C6848 XA6/XA3/MP0/a_216_n18# VREF 0.02fF
C6849 XA0/XA6/MP3/S VREF 0.02fF
C6850 XA7/XA1/XA5/MP1/S XA7/XA4/A 0.02fF
C6851 XA5/XA9/B XA5/XA9/MP1/a_216_334# 0.08fF
C6852 XB2/XA3/MP0/a_216_n18# AVDD 0.08fF
C6853 XA1/XA1/XA2/Y XA1/CN1 0.04fF
C6854 XA1/XA2/A XA1/XA2/MN3/a_324_n18# 0.15fF
C6855 XA7/XA1/XA5/MP2/a_216_n18# XA7/XA1/XA5/MP1/a_216_n18# 0.01fF
C6856 XA5/CP0 XA5/XA4/MP1/a_216_n18# 0.02fF
C6857 XDAC1/XC128b<2>/XRES2/B XDAC1/X16ab/XRES16/B 0.01fF
C6858 XA8/XA3/MP1/a_216_n18# XA8/XA3/MP0/a_216_n18# 0.01fF
C6859 XA3/XA1/XA1/MP3/S AVSS 0.02fF
C6860 XA6/XA1/XA1/MN1/a_324_n18# XA6/EN 0.08fF
C6861 XB1/XCAPB1/XCAPB1/m3_252_308# XB1/XA3/B 0.02fF
C6862 XA20/CPO XA2/XA1/XA1/MP2/a_216_n18# 0.06fF
C6863 XA8/XA5/MN2/a_324_n18# XA8/CP0 0.15fF
C6864 XA8/XA11/MP1/a_216_n18# AVDD 0.08fF
C6865 XA0/XA1/XA2/Y XA0/XA1/XA4/MN0/a_324_n18# 0.02fF
C6866 XA4/XA5/MN3/a_324_n18# XA4/XA6/MN0/a_324_n18# 0.01fF
C6867 XA2/XA4/MN1/a_324_n18# XA2/XA4/MN0/a_324_n18# 0.01fF
C6868 XB2/XA3/MP2/a_216_n18# XB2/CKN 0.07fF
C6869 XA4/CN0 SARP 0.02fF
C6870 XA5/XA6/MP0/a_216_n18# VREF 0.01fF
C6871 XA8/ENO XA8/XA9/B 0.07fF
C6872 XA2/XA2/A XA2/XA2/MP3/a_216_n18# 0.15fF
C6873 XA7/XA12/A AVDD 0.44fF
C6874 XA1/XA1/XA1/MP0/a_216_n18# XA1/EN 0.01fF
C6875 XA6/XA6/MP1/S CK_SAMPLE 0.03fF
C6876 XA2/CP0 XA2/XA4/MN2/a_324_n18# 0.01fF
C6877 VREF XA3/XA4/MP2/a_216_n18# 0.03fF
C6878 XA3/XA9/MN1/S AVSS 0.15fF
C6879 XA1/EN XA2/XA1/XA2/Y 0.02fF
C6880 XA3/CEO XA4/XA11/MN1/a_324_n18# 0.08fF
C6881 XA20/XA4/MN5/a_324_n18# XA20/XA4/MN6/a_324_n18# 0.01fF
C6882 XA20/CPO XA0/XA1/XA1/MP3/a_216_n18# 0.08fF
C6883 XA1/XA4/A XA2/CN1 0.07fF
C6884 XA8/XA1/XA1/MP2/S XA8/ENO 0.14fF
C6885 XA1/XA3/MP0/a_216_n18# AVDD 0.08fF
C6886 XA0/XA7/MN0/a_324_n18# XA0/XA9/B 0.01fF
C6887 XA5/CN0 SARP 0.02fF
C6888 XA0/XA1/XA4/MP1/a_216_n18# AVDD 0.08fF
C6889 XA4/XA2/MP3/a_216_n18# AVDD 0.07fF
C6890 XA2/EN XA2/CP0 0.02fF
C6891 D<1> XDAC1/XC32a<0>/XRES16/B 0.02fF
C6892 XA7/XA9/MP1/a_216_334# XA7/XA9/Y 0.07fF
C6893 XA20/XA3/MP6/a_216_n18# XA20/XA4/MP0/a_216_n18# 0.01fF
C6894 XA0/XA1/XA2/Y AVSS 0.27fF
C6895 XA4/EN AVDD 4.11fF
C6896 XA8/ENO XA8/XA6/MP3/S 0.02fF
C6897 XA2/XA7/MN0/a_324_n18# AVSS 0.01fF
C6898 XA8/XA7/MN0/a_324_n18# AVSS 0.01fF
C6899 XA2/XA3/MN1/a_324_n18# XA2/CN1 0.16fF
C6900 XA20/XA2/N2 XA20/CPO 0.12fF
C6901 XA4/XA5/MP2/a_216_n18# AVDD 0.07fF
C6902 XB1/XCAPB1/XCAPB0/m3_324_308# XB1/XA4/GNG 0.07fF
C6903 XA0/CP0 XA2/CN1 0.10fF
C6904 XB2/XCAPB1/XCAPB4/m3_9828_132# XB2/XA4/GNG 0.03fF
C6905 XA6/XA5/MN3/a_324_n18# XA6/CP0 0.15fF
C6906 XA6/XA2/A XA6/XA2/MN1/a_324_n18# 0.15fF
C6907 XA2/XA9/Y XA2/CEO 0.01fF
C6908 XA4/XA1/XA1/MP2/S AVDD 0.11fF
C6909 XA0/XA13/MN1/a_324_n18# AVSS 0.09fF
C6910 XA7/XA6/MN0/a_324_n18# AVSS 0.01fF
C6911 XA0/XA9/B XA0/CN0 0.07fF
C6912 XA6/XA1/XA1/MN3/a_324_n18# XA7/EN 0.01fF
C6913 XA2/XA13/MN1/a_324_334# AVSS 0.10fF
C6914 XA20/XA12/MN0/a_324_n18# XA20/XA11/MN1/a_324_n18# 0.01fF
C6915 XA3/CN0 XA0/CN0 0.11fF
C6916 XA6/CN0 XA6/XA5/MP3/a_216_n18# 0.02fF
C6917 SARN XB1/M4/G 0.17fF
C6918 XA1/XA1/XA1/MP2/a_216_n18# XA1/XA1/XA1/MP3/a_216_n18# 0.01fF
C6919 XA20/XA10/MP1/a_216_n18# XA20/XA9/MP0/a_216_334# 0.01fF
C6920 XA20/CNO XA2/XA1/XA1/MP1/a_216_n18# 0.06fF
C6921 XA4/XA6/MP1/S D<4> 0.02fF
C6922 XA2/CN0 AVDD 5.95fF
C6923 XA2/XA7/MN0/a_324_n18# XA2/XA9/B 0.01fF
C6924 XA3/XA2/A XA3/XA2/MN0/a_324_n18# 0.08fF
C6925 XA4/XA1/XA2/Y XA4/EN 0.14fF
C6926 XA0/XA2/A XA0/XA2/MP3/a_216_n18# 0.15fF
C6927 XA7/XA2/MN1/a_324_n18# XA7/XA2/A 0.15fF
C6928 XA8/CN0 XA8/XA9/B 0.07fF
C6929 XA7/XA11/A XA7/XA12/A 0.07fF
C6930 XA20/XA2/N2 XA20/XA3/N1 0.58fF
C6931 XA0/CP1 XDAC1/XC0/XRES16/B 0.22fF
C6932 XDAC2/X16ab/XRES1A/B AVSS 2.95fF
C6933 XA2/XA4/MP1/a_216_n18# VREF 0.02fF
C6934 XA3/EN XA2/XA1/XA5/MP1/S 0.02fF
C6935 XA2/XA9/MP1/a_216_n18# XA2/XA9/A 0.08fF
C6936 XDAC1/XC64a<0>/XRES8/B XDAC1/XC64a<0>/XRES1A/B 0.12fF
C6937 SAR_IP CK_SAMPLE_BSSW 0.04fF
C6938 XB2/M4/G XB2/XA4/MP1/a_216_n18# 0.08fF
C6939 XA4/XA3/MP2/a_216_n18# AVDD 0.07fF
C6940 D<8> XA1/CN1 0.69fF
C6941 XDAC2/XC64b<1>/XRES2/B SARN 3.05fF
C6942 XA0/CP0 XA0/XA6/MN0/a_324_n18# 0.07fF
C6943 XA7/XA6/MP3/S VREF 0.02fF
C6944 SARN XDAC2/XC32a<0>/XRES2/B 3.05fF
C6945 XA20/CPO XA20/XA3a/A 0.21fF
C6946 XA20/CNO XA0/XA1/XA1/MP1/a_216_n18# 0.06fF
C6947 XA6/XA1/XA5/MN2/S EN 0.02fF
C6948 XA5/XA4/MN3/a_324_n18# XA5/XA4/A 0.15fF
C6949 XA6/XA5/MP0/a_216_n18# XA6/XA4/MP3/a_216_n18# 0.01fF
C6950 XDAC2/XC128b<2>/XRES8/B XDAC2/XC128a<1>/XRES4/B 0.01fF
C6951 XA1/XA1/XA4/MN2/S XA1/XA1/XA4/MN1/S 0.04fF
C6952 XA4/XA9/MN1/a_324_334# XA4/XA11/MN0/a_324_n18# 0.01fF
C6953 XA1/CP0 XA1/XA5/MN2/a_324_n18# 0.15fF
C6954 XA7/CN1 VREF 0.76fF
C6955 XA7/XA1/XA5/MN1/S XA7/XA4/A 0.02fF
C6956 XA5/CP0 XA5/XA6/MN0/a_324_n18# 0.07fF
C6957 XA8/ENO VREF 0.97fF
C6958 D<5> XA3/XA1/XA1/MN2/S 0.01fF
C6959 XA8/ENO XA8/XA1/XA1/MN3/a_324_n18# 0.01fF
C6960 XB1/M8/a_324_334# XB1/M8/a_324_n18# 0.01fF
C6961 XA7/XA2/MP2/a_216_n18# XA7/XA2/A 0.15fF
C6962 XA2/XA4/A XA1/CN1 0.07fF
C6963 D<1> XA20/CPO 0.07fF
C6964 SARN AVDD 0.68fF
C6965 XA20/CNO XA3/XA1/XA2/Y 0.22fF
C6966 XA4/XA1/XA4/MP0/a_216_n18# AVDD 0.08fF
C6967 XA7/XA6/MP3/a_216_n18# AVDD 0.08fF
C6968 XA8/XA9/MP0/a_216_n18# XA8/XA8/MP0/a_216_n18# 0.01fF
C6969 XA0/XA4/A XA0/XA4/MP3/a_216_n18# 0.15fF
C6970 XA20/CPO XA0/XA1/XA2/MN0/a_324_n18# 0.01fF
C6971 XA1/CP0 XA1/XA5/MN0/a_324_n18# 0.09fF
C6972 XA5/XA6/MN1/S AVDD 0.01fF
C6973 XB1/XA2/MP0/G XB1/XA7/MN1/a_324_334# 0.07fF
C6974 XA0/XA1/XA2/MP0/a_216_n18# XA0/XA1/XA1/MP3/G 0.08fF
C6975 XA6/XA2/MN3/a_324_n18# XA6/XA2/A 0.15fF
C6976 XA20/XA3/N1 XA20/XA3a/A 0.29fF
C6977 XA3/XA2/A XA3/XA2/MN1/a_324_n18# 0.15fF
C6978 D<0> XA8/CP0 0.23fF
C6979 D<7> XA1/XA4/A 0.26fF
C6980 AVSS XB1/XA7/MN1/a_324_n18# 0.09fF
C6981 AVDD XA2/XA1/XA4/MN1/S 0.02fF
C6982 XA4/XA5/MP3/a_216_n18# XA4/CN0 0.02fF
C6983 XA8/EN XA8/XA1/XA5/MN2/a_324_n18# 0.08fF
C6984 XA20/XA2/MP3/a_216_n18# AVDD 0.18fF
C6985 XB1/XA5/MP1/a_216_n18# XB1/XA2/MP0/G 0.08fF
C6986 XB1/XA5b/MN1/a_324_n18# XB1/XA0/MN0/a_324_n18# 0.01fF
C6987 XA7/XA1/XA4/MP2/S XA7/XA4/A 0.05fF
C6988 XA20/XA2/MN2/a_324_n18# XA20/XA3/N1 0.01fF
C6989 XA2/XA2/A XA2/XA1/XA2/Y 0.01fF
C6990 XA2/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C6991 XA3/DONE XA3/XA9/B 0.03fF
C6992 XA8/XA7/MN0/a_324_n18# CK_SAMPLE 0.07fF
C6993 XA4/XA6/MP3/a_216_n18# AVDD 0.08fF
C6994 XA7/XA4/MN3/a_324_n18# XA7/CP0 0.02fF
C6995 XA8/XA9/MN1/S 0 0.05fF
C6996 XA8/XA9/MN1/a_324_n18# 0 0.15fF
C6997 XA8/XA9/Y 0 0.48fF
C6998 XA8/XA9/A 0 0.74fF
C6999 XA8/XA9/MP1/a_216_n18# 0 0.04fF
C7000 XA8/XA9/MN0/a_324_n18# 0 0.17fF
C7001 DONE 0 0.13fF
C7002 XA8/XA9/MP0/a_216_n18# 0 0.03fF
C7003 XA8/XA7/MN0/a_324_n18# 0 0.17fF
C7004 XA8/XA8/MN0/a_324_n18# 0 0.17fF
C7005 XA8/XA7/MP0/a_216_n18# 0 0.03fF
C7006 XA8/XA8/MP0/a_216_n18# 0 0.02fF
C7007 XA8/XA6/MN3/a_324_n18# 0 0.15fF
C7008 XA8/XA6/MN3/S 0 0.04fF
C7009 XA8/XA6/MN2/a_324_n18# 0 0.15fF
C7010 XA8/XA6/MN1/a_324_n18# 0 0.15fF
C7011 XA8/XA6/MP3/a_216_n18# 0 0.03fF
C7012 XA8/XA6/MN1/S 0 0.04fF
C7013 XA8/XA6/MN0/a_324_n18# 0 0.17fF
C7014 XA8/XA6/MP3/S 0 0.01fF
C7015 XA8/XA6/MP2/a_216_n18# 0 0.02fF
C7016 XA8/XA6/MP1/a_216_n18# 0 0.03fF
C7017 XA8/XA9/B 0 0.83fF
C7018 XA8/XA6/MP1/S 0 0.01fF
C7019 XA8/XA6/MP0/a_216_n18# 0 0.05fF
C7020 XA8/CP0 0 1.71fF
C7021 XA8/XA5/MN3/a_324_n18# 0 0.15fF
C7022 XA8/XA5/MN2/a_324_n18# 0 0.15fF
C7023 XA8/XA5/MN1/a_324_n18# 0 0.15fF
C7024 XA8/XA5/MP3/a_216_n18# 0 0.03fF
C7025 XA8/CN0 0 0.38fF
C7026 XA8/XA5/MP2/a_216_n18# 0 0.02fF
C7027 XA8/XA5/MP1/a_216_n18# 0 0.03fF
C7028 XA8/XA4/A 0 1.93fF
C7029 XA8/XA4/MN3/a_324_n18# 0 0.15fF
C7030 XA8/XA5/MN0/a_324_n18# 0 0.17fF
C7031 XA8/XA4/MN2/a_324_n18# 0 0.15fF
C7032 XA8/XA4/MN1/a_324_n18# 0 0.15fF
C7033 XA8/XA4/MP3/a_216_n18# 0 0.03fF
C7034 XA8/XA5/MP0/a_216_n18# 0 0.05fF
C7035 XA8/XA4/MP2/a_216_n18# 0 0.02fF
C7036 XA8/XA4/MP1/a_216_n18# 0 0.03fF
C7037 XA8/CN1 0 1.76fF
C7038 XA8/XA3/MN3/a_324_n18# 0 0.15fF
C7039 XA8/XA4/MN0/a_324_n18# 0 0.17fF
C7040 XA8/XA3/MN2/a_324_n18# 0 0.15fF
C7041 XA8/XA3/MN1/a_324_n18# 0 0.15fF
C7042 XA8/XA3/MP3/a_216_n18# 0 0.03fF
C7043 XA8/XA4/MP0/a_216_n18# 0 0.05fF
C7044 D<0> 0 0.35fF
C7045 XA8/XA3/MN0/a_324_n18# 0 0.17fF
C7046 XA8/XA3/MP2/a_216_n18# 0 0.02fF
C7047 XA8/XA3/MP1/a_216_n18# 0 0.03fF
C7048 XA8/XA3/MP0/a_216_n18# 0 0.05fF
C7049 XA8/XA2/A 0 1.31fF
C7050 XA8/XA2/MN3/a_324_n18# 0 0.15fF
C7051 XA8/XA2/MN2/a_324_n18# 0 0.15fF
C7052 XA8/XA2/MN1/a_324_n18# 0 0.15fF
C7053 XA8/XA2/MP3/a_216_n18# 0 0.03fF
C7054 XA8/XA2/MP2/a_216_n18# 0 0.02fF
C7055 XA8/XA2/MP1/a_216_n18# 0 0.03fF
C7056 XA8/XA1/XA5/MN2/S 0 0.06fF
C7057 XA8/XA2/MN0/a_324_n18# 0 0.17fF
C7058 XA8/XA1/XA5/MN1/S 0 0.06fF
C7059 XA8/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7060 XA8/XA1/XA5/MP2/S 0 0.02fF
C7061 XA8/XA2/MP0/a_216_n18# 0 0.05fF
C7062 XA8/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7063 XA8/XA1/XA5/MP1/S 0 0.02fF
C7064 XA8/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7065 XA8/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7066 XA8/XA1/XA4/MN2/S 0 0.06fF
C7067 XA8/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7068 XA8/XA1/XA4/MN1/S 0 0.06fF
C7069 XA8/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7070 XA8/XA1/XA4/MP2/S 0 0.02fF
C7071 XA8/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7072 XA8/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7073 XA8/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7074 XA8/XA1/XA4/MP1/S 0 0.02fF
C7075 XA8/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7076 XA8/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7077 XA8/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7078 XA8/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7079 XA8/XA1/XA2/Y 0 0.78fF
C7080 XA8/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7081 XA8/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7082 XA8/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7083 XA8/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7084 XA8/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7085 XA8/XA1/XA1/MP3/G 0 0.62fF
C7086 XA8/XA1/XA1/MN2/S 0 0.16fF
C7087 XA8/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7088 XA8/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7089 XA8/ENO 0 0.55fF
C7090 XA8/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7091 XA8/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7092 XA8/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7093 XA8/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7094 XA8/XA13/MN1/a_324_n18# 0 0.17fF
C7095 XA8/XA13/MN1/a_324_334# 0 0.32fF
C7096 XA8/XA13/MP1/a_216_n18# 0 0.03fF
C7097 XA8/XA13/MP1/a_216_334# 0 0.21fF
C7098 XA8/XA12/MN0/a_324_n18# 0 0.17fF
C7099 XA8/CEO 0 0.32fF
C7100 XA8/XA12/MP0/a_216_n18# 0 0.03fF
C7101 XA8/XA11/MN1/a_324_n18# 0 0.15fF
C7102 XA8/XA11/MP1/S 0 0.02fF
C7103 XA8/XA12/A 0 0.51fF
C7104 XA8/XA11/A 0 0.45fF
C7105 XA8/XA11/MP1/a_216_n18# 0 0.04fF
C7106 XA8/XA9/MN1/a_324_334# 0 0.17fF
C7107 XA8/XA11/MN0/a_324_n18# 0 0.17fF
C7108 XA8/XA9/MP1/a_216_334# 0 0.03fF
C7109 XA8/XA11/MP0/a_216_n18# 0 0.03fF
C7110 XA7/XA9/MN1/S 0 0.05fF
C7111 XA7/XA9/MN1/a_324_n18# 0 0.15fF
C7112 XA7/XA9/Y 0 0.48fF
C7113 XA7/XA9/A 0 0.74fF
C7114 XA7/XA9/MP1/a_216_n18# 0 0.04fF
C7115 XA7/XA9/MN0/a_324_n18# 0 0.17fF
C7116 XA7/DONE 0 0.07fF
C7117 XA7/XA9/MP0/a_216_n18# 0 0.03fF
C7118 XA7/XA7/MN0/a_324_n18# 0 0.17fF
C7119 XA7/XA8/MN0/a_324_n18# 0 0.17fF
C7120 XA7/XA7/MP0/a_216_n18# 0 0.03fF
C7121 XA7/XA8/MP0/a_216_n18# 0 0.02fF
C7122 XA7/XA6/MN3/a_324_n18# 0 0.15fF
C7123 XA7/XA6/MN3/S 0 0.04fF
C7124 XA7/XA6/MN2/a_324_n18# 0 0.15fF
C7125 XA7/XA6/MN1/a_324_n18# 0 0.15fF
C7126 XA7/XA6/MP3/a_216_n18# 0 0.03fF
C7127 XA7/XA6/MN1/S 0 0.04fF
C7128 XA7/XA6/MN0/a_324_n18# 0 0.17fF
C7129 XA7/XA6/MP3/S 0 0.01fF
C7130 XA7/XA6/MP2/a_216_n18# 0 0.02fF
C7131 XA7/XA6/MP1/a_216_n18# 0 0.03fF
C7132 XA7/XA9/B 0 0.83fF
C7133 XA7/XA6/MP1/S 0 0.01fF
C7134 XA7/XA6/MP0/a_216_n18# 0 0.05fF
C7135 XA7/CP0 0 1.71fF
C7136 XA7/XA5/MN3/a_324_n18# 0 0.15fF
C7137 XA7/XA5/MN2/a_324_n18# 0 0.15fF
C7138 XA7/XA5/MN1/a_324_n18# 0 0.15fF
C7139 XA7/XA5/MP3/a_216_n18# 0 0.03fF
C7140 XA7/CN0 0 5.50fF
C7141 XA7/XA5/MP2/a_216_n18# 0 0.02fF
C7142 XA7/XA5/MP1/a_216_n18# 0 0.03fF
C7143 XA7/XA4/A 0 1.93fF
C7144 XA7/XA4/MN3/a_324_n18# 0 0.15fF
C7145 XA7/XA5/MN0/a_324_n18# 0 0.17fF
C7146 XA7/XA4/MN2/a_324_n18# 0 0.15fF
C7147 XA7/XA4/MN1/a_324_n18# 0 0.15fF
C7148 XA7/XA4/MP3/a_216_n18# 0 0.03fF
C7149 XA7/XA5/MP0/a_216_n18# 0 0.05fF
C7150 XA7/XA4/MP2/a_216_n18# 0 0.02fF
C7151 XA7/XA4/MP1/a_216_n18# 0 0.03fF
C7152 XA7/CN1 0 1.76fF
C7153 XA7/XA3/MN3/a_324_n18# 0 0.15fF
C7154 XA7/XA4/MN0/a_324_n18# 0 0.17fF
C7155 XA7/XA3/MN2/a_324_n18# 0 0.15fF
C7156 XA7/XA3/MN1/a_324_n18# 0 0.15fF
C7157 XA7/XA3/MP3/a_216_n18# 0 0.03fF
C7158 XA7/XA4/MP0/a_216_n18# 0 0.05fF
C7159 D<1> 0 4.86fF
C7160 XA7/XA3/MN0/a_324_n18# 0 0.17fF
C7161 XA7/XA3/MP2/a_216_n18# 0 0.02fF
C7162 XA7/XA3/MP1/a_216_n18# 0 0.03fF
C7163 XA7/XA3/MP0/a_216_n18# 0 0.05fF
C7164 XA7/XA2/A 0 1.31fF
C7165 XA7/XA2/MN3/a_324_n18# 0 0.15fF
C7166 XA7/XA2/MN2/a_324_n18# 0 0.15fF
C7167 XA7/XA2/MN1/a_324_n18# 0 0.15fF
C7168 XA7/XA2/MP3/a_216_n18# 0 0.03fF
C7169 XA7/XA2/MP2/a_216_n18# 0 0.02fF
C7170 XA7/XA2/MP1/a_216_n18# 0 0.03fF
C7171 XA7/XA1/XA5/MN2/S 0 0.06fF
C7172 XA7/XA2/MN0/a_324_n18# 0 0.17fF
C7173 XA7/XA1/XA5/MN1/S 0 0.06fF
C7174 XA7/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7175 XA7/XA1/XA5/MP2/S 0 0.02fF
C7176 XA7/XA2/MP0/a_216_n18# 0 0.05fF
C7177 XA7/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7178 XA7/XA1/XA5/MP1/S 0 0.02fF
C7179 XA7/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7180 XA7/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7181 XA7/XA1/XA4/MN2/S 0 0.06fF
C7182 XA7/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7183 XA7/XA1/XA4/MN1/S 0 0.06fF
C7184 XA7/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7185 XA7/XA1/XA4/MP2/S 0 0.02fF
C7186 XA7/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7187 XA7/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7188 XA7/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7189 XA7/XA1/XA4/MP1/S 0 0.02fF
C7190 XA7/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7191 XA7/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7192 XA7/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7193 XA7/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7194 XA7/XA1/XA2/Y 0 0.78fF
C7195 XA7/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7196 XA7/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7197 XA7/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7198 XA7/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7199 XA7/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7200 XA7/XA1/XA1/MP3/G 0 0.62fF
C7201 XA7/XA1/XA1/MN2/S 0 0.16fF
C7202 XA7/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7203 XA7/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7204 XA8/EN 0 2.22fF
C7205 XA7/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7206 XA7/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7207 XA7/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7208 XA7/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7209 XA7/XA13/MN1/a_324_n18# 0 0.17fF
C7210 XA7/XA13/MN1/a_324_334# 0 0.32fF
C7211 XA7/XA13/MP1/a_216_n18# 0 0.03fF
C7212 XA7/XA13/MP1/a_216_334# 0 0.21fF
C7213 XA7/XA12/MN0/a_324_n18# 0 0.17fF
C7214 XA7/CEO 0 0.61fF
C7215 XA7/XA12/MP0/a_216_n18# 0 0.03fF
C7216 XA7/XA11/MN1/a_324_n18# 0 0.15fF
C7217 XA7/XA11/MP1/S 0 0.02fF
C7218 XA7/XA12/A 0 0.51fF
C7219 XA7/XA11/A 0 0.45fF
C7220 XA7/XA11/MP1/a_216_n18# 0 0.04fF
C7221 XA7/XA9/MN1/a_324_334# 0 0.17fF
C7222 XA7/XA11/MN0/a_324_n18# 0 0.17fF
C7223 XA7/XA9/MP1/a_216_334# 0 0.03fF
C7224 XA7/XA11/MP0/a_216_n18# 0 0.03fF
C7225 XA6/XA9/MN1/S 0 0.05fF
C7226 XA6/XA9/MN1/a_324_n18# 0 0.15fF
C7227 XA6/XA9/Y 0 0.48fF
C7228 XA6/XA9/A 0 0.74fF
C7229 XA6/XA9/MP1/a_216_n18# 0 0.04fF
C7230 XA6/XA9/MN0/a_324_n18# 0 0.17fF
C7231 XA6/DONE 0 0.07fF
C7232 XA6/XA9/MP0/a_216_n18# 0 0.03fF
C7233 XA6/XA7/MN0/a_324_n18# 0 0.17fF
C7234 XA6/XA8/MN0/a_324_n18# 0 0.17fF
C7235 XA6/XA7/MP0/a_216_n18# 0 0.03fF
C7236 XA6/XA8/MP0/a_216_n18# 0 0.02fF
C7237 XA6/XA6/MN3/a_324_n18# 0 0.15fF
C7238 XA6/XA6/MN3/S 0 0.04fF
C7239 XA6/XA6/MN2/a_324_n18# 0 0.15fF
C7240 XA6/XA6/MN1/a_324_n18# 0 0.15fF
C7241 XA6/XA6/MP3/a_216_n18# 0 0.03fF
C7242 XA6/XA6/MN1/S 0 0.04fF
C7243 XA6/XA6/MN0/a_324_n18# 0 0.17fF
C7244 XA6/XA6/MP3/S 0 0.01fF
C7245 XA6/XA6/MP2/a_216_n18# 0 0.02fF
C7246 XA6/XA6/MP1/a_216_n18# 0 0.03fF
C7247 XA6/XA9/B 0 0.83fF
C7248 XA6/XA6/MP1/S 0 0.01fF
C7249 XA6/XA6/MP0/a_216_n18# 0 0.05fF
C7250 XA6/CP0 0 1.71fF
C7251 XA6/XA5/MN3/a_324_n18# 0 0.15fF
C7252 XA6/XA5/MN2/a_324_n18# 0 0.15fF
C7253 XA6/XA5/MN1/a_324_n18# 0 0.15fF
C7254 XA6/XA5/MP3/a_216_n18# 0 0.03fF
C7255 XA6/CN0 0 3.04fF
C7256 XA6/XA5/MP2/a_216_n18# 0 0.02fF
C7257 XA6/XA5/MP1/a_216_n18# 0 0.03fF
C7258 XA6/XA4/A 0 1.93fF
C7259 XA6/XA4/MN3/a_324_n18# 0 0.15fF
C7260 XA6/XA5/MN0/a_324_n18# 0 0.17fF
C7261 XA6/XA4/MN2/a_324_n18# 0 0.15fF
C7262 XA6/XA4/MN1/a_324_n18# 0 0.15fF
C7263 XA6/XA4/MP3/a_216_n18# 0 0.03fF
C7264 XA6/XA5/MP0/a_216_n18# 0 0.05fF
C7265 XA6/XA4/MP2/a_216_n18# 0 0.02fF
C7266 XA6/XA4/MP1/a_216_n18# 0 0.03fF
C7267 XA6/CN1 0 1.76fF
C7268 XA6/XA3/MN3/a_324_n18# 0 0.15fF
C7269 XA6/XA4/MN0/a_324_n18# 0 0.17fF
C7270 XA6/XA3/MN2/a_324_n18# 0 0.15fF
C7271 XA6/XA3/MN1/a_324_n18# 0 0.15fF
C7272 XA6/XA3/MP3/a_216_n18# 0 0.03fF
C7273 XA6/XA4/MP0/a_216_n18# 0 0.05fF
C7274 D<2> 0 4.37fF
C7275 XA6/XA3/MN0/a_324_n18# 0 0.17fF
C7276 XA6/XA3/MP2/a_216_n18# 0 0.02fF
C7277 XA6/XA3/MP1/a_216_n18# 0 0.03fF
C7278 XA6/XA3/MP0/a_216_n18# 0 0.05fF
C7279 XA6/XA2/A 0 1.31fF
C7280 XA6/XA2/MN3/a_324_n18# 0 0.15fF
C7281 XA6/XA2/MN2/a_324_n18# 0 0.15fF
C7282 XA6/XA2/MN1/a_324_n18# 0 0.15fF
C7283 XA6/XA2/MP3/a_216_n18# 0 0.03fF
C7284 XA6/XA2/MP2/a_216_n18# 0 0.02fF
C7285 XA6/XA2/MP1/a_216_n18# 0 0.03fF
C7286 XA6/XA1/XA5/MN2/S 0 0.06fF
C7287 XA6/XA2/MN0/a_324_n18# 0 0.17fF
C7288 XA6/XA1/XA5/MN1/S 0 0.06fF
C7289 XA6/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7290 XA6/XA1/XA5/MP2/S 0 0.02fF
C7291 XA6/XA2/MP0/a_216_n18# 0 0.05fF
C7292 XA6/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7293 XA6/XA1/XA5/MP1/S 0 0.02fF
C7294 XA6/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7295 XA6/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7296 XA6/XA1/XA4/MN2/S 0 0.06fF
C7297 XA6/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7298 XA6/XA1/XA4/MN1/S 0 0.06fF
C7299 XA6/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7300 XA6/XA1/XA4/MP2/S 0 0.02fF
C7301 XA6/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7302 XA6/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7303 XA6/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7304 XA6/XA1/XA4/MP1/S 0 0.02fF
C7305 XA6/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7306 XA6/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7307 XA6/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7308 XA6/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7309 XA6/XA1/XA2/Y 0 0.78fF
C7310 XA6/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7311 XA6/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7312 XA6/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7313 XA6/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7314 XA6/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7315 XA6/XA1/XA1/MP3/G 0 0.62fF
C7316 XA6/XA1/XA1/MN2/S 0 0.16fF
C7317 XA6/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7318 XA6/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7319 XA7/EN 0 2.02fF
C7320 XA6/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7321 XA6/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7322 XA6/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7323 XA6/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7324 XA6/XA13/MN1/a_324_n18# 0 0.17fF
C7325 XA6/XA13/MN1/a_324_334# 0 0.32fF
C7326 XA6/XA13/MP1/a_216_n18# 0 0.03fF
C7327 XA6/XA13/MP1/a_216_334# 0 0.21fF
C7328 XA6/XA12/MN0/a_324_n18# 0 0.17fF
C7329 XA6/CEO 0 0.42fF
C7330 XA6/XA12/MP0/a_216_n18# 0 0.03fF
C7331 XA6/XA11/MN1/a_324_n18# 0 0.15fF
C7332 XA6/XA11/MP1/S 0 0.02fF
C7333 XA6/XA12/A 0 0.51fF
C7334 XA6/XA11/A 0 0.45fF
C7335 XA6/XA11/MP1/a_216_n18# 0 0.04fF
C7336 XA6/XA9/MN1/a_324_334# 0 0.17fF
C7337 XA6/XA11/MN0/a_324_n18# 0 0.17fF
C7338 XA6/XA9/MP1/a_216_334# 0 0.03fF
C7339 XA6/XA11/MP0/a_216_n18# 0 0.03fF
C7340 XA5/XA9/MN1/S 0 0.05fF
C7341 XA5/XA9/MN1/a_324_n18# 0 0.15fF
C7342 XA5/XA9/Y 0 0.48fF
C7343 XA5/XA9/A 0 0.74fF
C7344 XA5/XA9/MP1/a_216_n18# 0 0.04fF
C7345 XA5/XA9/MN0/a_324_n18# 0 0.17fF
C7346 XA5/DONE 0 0.07fF
C7347 XA5/XA9/MP0/a_216_n18# 0 0.03fF
C7348 XA5/XA7/MN0/a_324_n18# 0 0.17fF
C7349 XA5/XA8/MN0/a_324_n18# 0 0.17fF
C7350 XA5/XA7/MP0/a_216_n18# 0 0.03fF
C7351 XA5/XA8/MP0/a_216_n18# 0 0.02fF
C7352 XA5/XA6/MN3/a_324_n18# 0 0.15fF
C7353 XA5/XA6/MN3/S 0 0.04fF
C7354 XA5/XA6/MN2/a_324_n18# 0 0.15fF
C7355 XA5/XA6/MN1/a_324_n18# 0 0.15fF
C7356 XA5/XA6/MP3/a_216_n18# 0 0.03fF
C7357 XA5/XA6/MN1/S 0 0.04fF
C7358 XA5/XA6/MN0/a_324_n18# 0 0.17fF
C7359 XA5/XA6/MP3/S 0 0.01fF
C7360 XA5/XA6/MP2/a_216_n18# 0 0.02fF
C7361 XA5/XA6/MP1/a_216_n18# 0 0.03fF
C7362 XA5/XA9/B 0 0.83fF
C7363 XA5/XA6/MP1/S 0 0.01fF
C7364 XA5/XA6/MP0/a_216_n18# 0 0.05fF
C7365 XA5/CP0 0 1.71fF
C7366 XA5/XA5/MN3/a_324_n18# 0 0.15fF
C7367 XA5/XA5/MN2/a_324_n18# 0 0.15fF
C7368 XA5/XA5/MN1/a_324_n18# 0 0.15fF
C7369 XA5/XA5/MP3/a_216_n18# 0 0.03fF
C7370 XA5/CN0 0 2.23fF
C7371 XA5/XA5/MP2/a_216_n18# 0 0.02fF
C7372 XA5/XA5/MP1/a_216_n18# 0 0.03fF
C7373 XA5/XA4/A 0 1.93fF
C7374 XA5/XA4/MN3/a_324_n18# 0 0.15fF
C7375 XA5/XA5/MN0/a_324_n18# 0 0.17fF
C7376 XA5/XA4/MN2/a_324_n18# 0 0.15fF
C7377 XA5/XA4/MN1/a_324_n18# 0 0.15fF
C7378 XA5/XA4/MP3/a_216_n18# 0 0.03fF
C7379 XA5/XA5/MP0/a_216_n18# 0 0.05fF
C7380 XA5/XA4/MP2/a_216_n18# 0 0.02fF
C7381 XA5/XA4/MP1/a_216_n18# 0 0.03fF
C7382 XA5/CN1 0 1.76fF
C7383 XA5/XA3/MN3/a_324_n18# 0 0.15fF
C7384 XA5/XA4/MN0/a_324_n18# 0 0.17fF
C7385 XA5/XA3/MN2/a_324_n18# 0 0.15fF
C7386 XA5/XA3/MN1/a_324_n18# 0 0.15fF
C7387 XA5/XA3/MP3/a_216_n18# 0 0.03fF
C7388 XA5/XA4/MP0/a_216_n18# 0 0.05fF
C7389 D<3> 0 2.63fF
C7390 XA5/XA3/MN0/a_324_n18# 0 0.17fF
C7391 XA5/XA3/MP2/a_216_n18# 0 0.02fF
C7392 XA5/XA3/MP1/a_216_n18# 0 0.03fF
C7393 XA5/XA3/MP0/a_216_n18# 0 0.05fF
C7394 XA5/XA2/A 0 1.31fF
C7395 XA5/XA2/MN3/a_324_n18# 0 0.15fF
C7396 XA5/XA2/MN2/a_324_n18# 0 0.15fF
C7397 XA5/XA2/MN1/a_324_n18# 0 0.15fF
C7398 XA5/XA2/MP3/a_216_n18# 0 0.03fF
C7399 XA5/XA2/MP2/a_216_n18# 0 0.02fF
C7400 XA5/XA2/MP1/a_216_n18# 0 0.03fF
C7401 XA5/XA1/XA5/MN2/S 0 0.06fF
C7402 XA5/XA2/MN0/a_324_n18# 0 0.17fF
C7403 XA5/XA1/XA5/MN1/S 0 0.06fF
C7404 XA5/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7405 XA5/XA1/XA5/MP2/S 0 0.02fF
C7406 XA5/XA2/MP0/a_216_n18# 0 0.05fF
C7407 XA5/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7408 XA5/XA1/XA5/MP1/S 0 0.02fF
C7409 XA5/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7410 XA5/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7411 XA5/XA1/XA4/MN2/S 0 0.06fF
C7412 XA5/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7413 XA5/XA1/XA4/MN1/S 0 0.06fF
C7414 XA5/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7415 XA5/XA1/XA4/MP2/S 0 0.02fF
C7416 XA5/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7417 XA5/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7418 XA5/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7419 XA5/XA1/XA4/MP1/S 0 0.02fF
C7420 XA5/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7421 XA5/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7422 XA5/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7423 XA5/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7424 XA5/XA1/XA2/Y 0 0.78fF
C7425 XA5/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7426 XA5/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7427 XA5/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7428 XA5/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7429 XA5/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7430 XA5/XA1/XA1/MP3/G 0 0.62fF
C7431 XA5/XA1/XA1/MN2/S 0 0.16fF
C7432 XA5/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7433 XA5/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7434 XA6/EN 0 2.11fF
C7435 XA5/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7436 XA5/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7437 XA5/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7438 XA5/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7439 XA5/XA13/MN1/a_324_n18# 0 0.17fF
C7440 XA5/XA13/MN1/a_324_334# 0 0.32fF
C7441 XA5/XA13/MP1/a_216_n18# 0 0.03fF
C7442 XA5/XA13/MP1/a_216_334# 0 0.21fF
C7443 XA5/XA12/MN0/a_324_n18# 0 0.17fF
C7444 XA5/CEO 0 0.61fF
C7445 XA5/XA12/MP0/a_216_n18# 0 0.03fF
C7446 XA5/XA11/MN1/a_324_n18# 0 0.15fF
C7447 XA5/XA11/MP1/S 0 0.02fF
C7448 XA5/XA12/A 0 0.51fF
C7449 XA5/XA11/A 0 0.45fF
C7450 XA5/XA11/MP1/a_216_n18# 0 0.04fF
C7451 XA5/XA9/MN1/a_324_334# 0 0.17fF
C7452 XA5/XA11/MN0/a_324_n18# 0 0.17fF
C7453 XA5/XA9/MP1/a_216_334# 0 0.03fF
C7454 XA5/XA11/MP0/a_216_n18# 0 0.03fF
C7455 XA4/XA9/MN1/S 0 0.05fF
C7456 XA4/XA9/MN1/a_324_n18# 0 0.15fF
C7457 XA4/XA9/Y 0 0.48fF
C7458 XA4/XA9/A 0 0.74fF
C7459 XA4/XA9/MP1/a_216_n18# 0 0.04fF
C7460 XA4/XA9/MN0/a_324_n18# 0 0.17fF
C7461 XA4/DONE 0 0.07fF
C7462 XA4/XA9/MP0/a_216_n18# 0 0.03fF
C7463 XA4/XA7/MN0/a_324_n18# 0 0.17fF
C7464 XA4/XA8/MN0/a_324_n18# 0 0.17fF
C7465 XA4/XA7/MP0/a_216_n18# 0 0.03fF
C7466 XA4/XA8/MP0/a_216_n18# 0 0.02fF
C7467 XA4/XA6/MN3/a_324_n18# 0 0.15fF
C7468 XA4/XA6/MN3/S 0 0.04fF
C7469 XA4/XA6/MN2/a_324_n18# 0 0.15fF
C7470 XA4/XA6/MN1/a_324_n18# 0 0.15fF
C7471 XA4/XA6/MP3/a_216_n18# 0 0.03fF
C7472 XA4/XA6/MN1/S 0 0.04fF
C7473 XA4/XA6/MN0/a_324_n18# 0 0.17fF
C7474 XA4/XA6/MP3/S 0 0.01fF
C7475 XA4/XA6/MP2/a_216_n18# 0 0.02fF
C7476 XA4/XA6/MP1/a_216_n18# 0 0.03fF
C7477 XA4/XA9/B 0 0.83fF
C7478 XA4/XA6/MP1/S 0 0.01fF
C7479 XA4/XA6/MP0/a_216_n18# 0 0.05fF
C7480 XA4/CP0 0 1.71fF
C7481 XA4/XA5/MN3/a_324_n18# 0 0.15fF
C7482 XA4/XA5/MN2/a_324_n18# 0 0.15fF
C7483 XA4/XA5/MN1/a_324_n18# 0 0.15fF
C7484 XA4/XA5/MP3/a_216_n18# 0 0.03fF
C7485 XA4/CN0 0 3.02fF
C7486 XA4/XA5/MP2/a_216_n18# 0 0.02fF
C7487 XA4/XA5/MP1/a_216_n18# 0 0.03fF
C7488 XA4/XA4/A 0 1.93fF
C7489 XA4/XA4/MN3/a_324_n18# 0 0.15fF
C7490 XA4/XA5/MN0/a_324_n18# 0 0.17fF
C7491 XA4/XA4/MN2/a_324_n18# 0 0.15fF
C7492 XA4/XA4/MN1/a_324_n18# 0 0.15fF
C7493 XA4/XA4/MP3/a_216_n18# 0 0.03fF
C7494 XA4/XA5/MP0/a_216_n18# 0 0.05fF
C7495 XA4/XA4/MP2/a_216_n18# 0 0.02fF
C7496 XA4/XA4/MP1/a_216_n18# 0 0.03fF
C7497 XA4/CN1 0 1.76fF
C7498 XA4/XA3/MN3/a_324_n18# 0 0.15fF
C7499 XA4/XA4/MN0/a_324_n18# 0 0.17fF
C7500 XA4/XA3/MN2/a_324_n18# 0 0.15fF
C7501 XA4/XA3/MN1/a_324_n18# 0 0.15fF
C7502 XA4/XA3/MP3/a_216_n18# 0 0.03fF
C7503 XA4/XA4/MP0/a_216_n18# 0 0.05fF
C7504 D<4> 0 3.25fF
C7505 XA4/XA3/MN0/a_324_n18# 0 0.17fF
C7506 XA4/XA3/MP2/a_216_n18# 0 0.02fF
C7507 XA4/XA3/MP1/a_216_n18# 0 0.03fF
C7508 XA4/XA3/MP0/a_216_n18# 0 0.05fF
C7509 XA4/XA2/A 0 1.31fF
C7510 XA4/XA2/MN3/a_324_n18# 0 0.15fF
C7511 XA4/XA2/MN2/a_324_n18# 0 0.15fF
C7512 XA4/XA2/MN1/a_324_n18# 0 0.15fF
C7513 XA4/XA2/MP3/a_216_n18# 0 0.03fF
C7514 XA4/XA2/MP2/a_216_n18# 0 0.02fF
C7515 XA4/XA2/MP1/a_216_n18# 0 0.03fF
C7516 XA4/XA1/XA5/MN2/S 0 0.06fF
C7517 XA4/XA2/MN0/a_324_n18# 0 0.17fF
C7518 XA4/XA1/XA5/MN1/S 0 0.06fF
C7519 XA4/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7520 XA4/XA1/XA5/MP2/S 0 0.02fF
C7521 XA4/XA2/MP0/a_216_n18# 0 0.05fF
C7522 XA4/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7523 XA4/XA1/XA5/MP1/S 0 0.02fF
C7524 XA4/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7525 XA4/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7526 XA4/XA1/XA4/MN2/S 0 0.06fF
C7527 XA4/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7528 XA4/XA1/XA4/MN1/S 0 0.06fF
C7529 XA4/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7530 XA4/XA1/XA4/MP2/S 0 0.02fF
C7531 XA4/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7532 XA4/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7533 XA4/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7534 XA4/XA1/XA4/MP1/S 0 0.02fF
C7535 XA4/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7536 XA4/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7537 XA4/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7538 XA4/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7539 XA4/XA1/XA2/Y 0 0.78fF
C7540 XA4/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7541 XA4/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7542 XA4/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7543 XA4/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7544 XA4/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7545 XA4/XA1/XA1/MP3/G 0 0.62fF
C7546 XA4/XA1/XA1/MN2/S 0 0.16fF
C7547 XA4/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7548 XA4/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7549 XA5/EN 0 2.21fF
C7550 XA4/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7551 XA4/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7552 XA4/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7553 XA4/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7554 XA4/XA13/MN1/a_324_n18# 0 0.17fF
C7555 XA4/XA13/MN1/a_324_334# 0 0.32fF
C7556 XA4/XA13/MP1/a_216_n18# 0 0.03fF
C7557 XA4/XA13/MP1/a_216_334# 0 0.21fF
C7558 XA4/XA12/MN0/a_324_n18# 0 0.17fF
C7559 XA4/CEO 0 0.40fF
C7560 XA4/XA12/MP0/a_216_n18# 0 0.03fF
C7561 XA4/XA11/MN1/a_324_n18# 0 0.15fF
C7562 XA4/XA11/MP1/S 0 0.02fF
C7563 XA4/XA12/A 0 0.51fF
C7564 XA4/XA11/A 0 0.45fF
C7565 XA4/XA11/MP1/a_216_n18# 0 0.04fF
C7566 XA4/XA9/MN1/a_324_334# 0 0.17fF
C7567 XA4/XA11/MN0/a_324_n18# 0 0.17fF
C7568 XA4/XA9/MP1/a_216_334# 0 0.03fF
C7569 XA4/XA11/MP0/a_216_n18# 0 0.03fF
C7570 XA3/XA9/MN1/S 0 0.05fF
C7571 XA3/XA9/MN1/a_324_n18# 0 0.15fF
C7572 XA3/XA9/Y 0 0.48fF
C7573 XA3/XA9/A 0 0.74fF
C7574 XA3/XA9/MP1/a_216_n18# 0 0.04fF
C7575 XA3/XA9/MN0/a_324_n18# 0 0.17fF
C7576 XA3/DONE 0 0.07fF
C7577 XA3/XA9/MP0/a_216_n18# 0 0.03fF
C7578 XA3/XA7/MN0/a_324_n18# 0 0.17fF
C7579 XA3/XA8/MN0/a_324_n18# 0 0.17fF
C7580 XA3/XA7/MP0/a_216_n18# 0 0.03fF
C7581 XA3/XA8/MP0/a_216_n18# 0 0.02fF
C7582 XA3/XA6/MN3/a_324_n18# 0 0.15fF
C7583 XA3/XA6/MN3/S 0 0.04fF
C7584 XA3/XA6/MN2/a_324_n18# 0 0.15fF
C7585 XA3/XA6/MN1/a_324_n18# 0 0.15fF
C7586 XA3/XA6/MP3/a_216_n18# 0 0.03fF
C7587 XA3/XA6/MN1/S 0 0.04fF
C7588 XA3/XA6/MN0/a_324_n18# 0 0.17fF
C7589 XA3/XA6/MP3/S 0 0.01fF
C7590 XA3/XA6/MP2/a_216_n18# 0 0.02fF
C7591 XA3/XA6/MP1/a_216_n18# 0 0.03fF
C7592 XA3/XA9/B 0 0.83fF
C7593 XA3/XA6/MP1/S 0 0.01fF
C7594 XA3/XA6/MP0/a_216_n18# 0 0.05fF
C7595 XA3/CP0 0 4.28fF
C7596 XA3/XA5/MN3/a_324_n18# 0 0.15fF
C7597 XA3/XA5/MN2/a_324_n18# 0 0.15fF
C7598 XA3/XA5/MN1/a_324_n18# 0 0.15fF
C7599 XA3/XA5/MP3/a_216_n18# 0 0.03fF
C7600 XA3/CN0 0 2.90fF
C7601 XA3/XA5/MP2/a_216_n18# 0 0.02fF
C7602 XA3/XA5/MP1/a_216_n18# 0 0.03fF
C7603 XA3/XA4/A 0 1.93fF
C7604 XA3/XA4/MN3/a_324_n18# 0 0.15fF
C7605 XA3/XA5/MN0/a_324_n18# 0 0.17fF
C7606 XA3/XA4/MN2/a_324_n18# 0 0.15fF
C7607 XA3/XA4/MN1/a_324_n18# 0 0.15fF
C7608 XA3/XA4/MP3/a_216_n18# 0 0.03fF
C7609 XA3/XA5/MP0/a_216_n18# 0 0.05fF
C7610 XA3/XA4/MP2/a_216_n18# 0 0.02fF
C7611 XA3/XA4/MP1/a_216_n18# 0 0.03fF
C7612 XA3/XA3/MN3/a_324_n18# 0 0.15fF
C7613 XA3/XA4/MN0/a_324_n18# 0 0.17fF
C7614 XA3/XA3/MN2/a_324_n18# 0 0.15fF
C7615 XA3/XA3/MN1/a_324_n18# 0 0.15fF
C7616 XA3/XA3/MP3/a_216_n18# 0 0.03fF
C7617 XA3/XA4/MP0/a_216_n18# 0 0.05fF
C7618 XA3/XA3/MN0/a_324_n18# 0 0.17fF
C7619 XA3/XA3/MP2/a_216_n18# 0 0.02fF
C7620 XA3/XA3/MP1/a_216_n18# 0 0.03fF
C7621 XA3/XA3/MP0/a_216_n18# 0 0.05fF
C7622 XA3/XA2/A 0 1.31fF
C7623 XA3/XA2/MN3/a_324_n18# 0 0.15fF
C7624 XA3/XA2/MN2/a_324_n18# 0 0.15fF
C7625 XA3/XA2/MN1/a_324_n18# 0 0.15fF
C7626 XA3/XA2/MP3/a_216_n18# 0 0.03fF
C7627 XA3/XA2/MP2/a_216_n18# 0 0.02fF
C7628 XA3/XA2/MP1/a_216_n18# 0 0.03fF
C7629 XA3/XA1/XA5/MN2/S 0 0.06fF
C7630 XA3/XA2/MN0/a_324_n18# 0 0.17fF
C7631 XA3/XA1/XA5/MN1/S 0 0.06fF
C7632 XA3/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7633 XA3/XA1/XA5/MP2/S 0 0.02fF
C7634 XA3/XA2/MP0/a_216_n18# 0 0.05fF
C7635 XA3/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7636 XA3/XA1/XA5/MP1/S 0 0.02fF
C7637 XA3/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7638 XA3/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7639 XA3/XA1/XA4/MN2/S 0 0.06fF
C7640 XA3/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7641 XA3/XA1/XA4/MN1/S 0 0.06fF
C7642 XA3/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7643 XA3/XA1/XA4/MP2/S 0 0.02fF
C7644 XA3/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7645 XA3/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7646 XA3/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7647 XA3/XA1/XA4/MP1/S 0 0.02fF
C7648 XA3/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7649 XA3/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7650 XA3/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7651 XA3/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7652 XA3/XA1/XA2/Y 0 0.78fF
C7653 XA3/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7654 XA3/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7655 XA3/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7656 XA3/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7657 XA3/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7658 XA3/XA1/XA1/MP3/G 0 0.62fF
C7659 XA3/XA1/XA1/MN2/S 0 0.16fF
C7660 XA3/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7661 XA3/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7662 XA4/EN 0 2.27fF
C7663 XA3/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7664 XA3/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7665 XA3/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7666 XA3/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7667 XA3/XA13/MN1/a_324_n18# 0 0.17fF
C7668 XA3/XA13/MN1/a_324_334# 0 0.32fF
C7669 XA3/XA13/MP1/a_216_n18# 0 0.03fF
C7670 XA3/XA13/MP1/a_216_334# 0 0.21fF
C7671 XA3/XA12/MN0/a_324_n18# 0 0.17fF
C7672 XA3/CEO 0 0.55fF
C7673 XA3/XA12/MP0/a_216_n18# 0 0.03fF
C7674 XA3/XA11/MN1/a_324_n18# 0 0.15fF
C7675 XA3/XA11/MP1/S 0 0.02fF
C7676 XA3/XA12/A 0 0.51fF
C7677 XA3/XA11/A 0 0.45fF
C7678 XA3/XA11/MP1/a_216_n18# 0 0.04fF
C7679 XA3/XA9/MN1/a_324_334# 0 0.17fF
C7680 XA3/XA11/MN0/a_324_n18# 0 0.17fF
C7681 XA3/XA9/MP1/a_216_334# 0 0.03fF
C7682 XA3/XA11/MP0/a_216_n18# 0 0.03fF
C7683 XA2/XA9/MN1/S 0 0.05fF
C7684 XA2/XA9/MN1/a_324_n18# 0 0.15fF
C7685 XA2/XA9/Y 0 0.48fF
C7686 XA2/XA9/A 0 0.74fF
C7687 XA2/XA9/MP1/a_216_n18# 0 0.04fF
C7688 XA2/XA9/MN0/a_324_n18# 0 0.17fF
C7689 XA2/DONE 0 0.07fF
C7690 XA2/XA9/MP0/a_216_n18# 0 0.03fF
C7691 XA2/XA7/MN0/a_324_n18# 0 0.17fF
C7692 XA2/XA8/MN0/a_324_n18# 0 0.17fF
C7693 XA2/XA7/MP0/a_216_n18# 0 0.03fF
C7694 XA2/XA8/MP0/a_216_n18# 0 0.02fF
C7695 XA2/XA6/MN3/a_324_n18# 0 0.15fF
C7696 XA2/XA6/MN3/S 0 0.04fF
C7697 XA2/XA6/MN2/a_324_n18# 0 0.15fF
C7698 XA2/XA6/MN1/a_324_n18# 0 0.15fF
C7699 XA2/XA6/MP3/a_216_n18# 0 0.03fF
C7700 XA2/XA6/MN1/S 0 0.04fF
C7701 XA2/XA6/MN0/a_324_n18# 0 0.17fF
C7702 XA2/XA6/MP3/S 0 0.01fF
C7703 XA2/XA6/MP2/a_216_n18# 0 0.02fF
C7704 XA2/XA6/MP1/a_216_n18# 0 0.03fF
C7705 XA2/XA9/B 0 0.83fF
C7706 XA2/XA6/MP1/S 0 0.01fF
C7707 XA2/XA6/MP0/a_216_n18# 0 0.05fF
C7708 XA2/CP0 0 4.37fF
C7709 XA2/XA5/MN3/a_324_n18# 0 0.15fF
C7710 XA2/XA5/MN2/a_324_n18# 0 0.15fF
C7711 XA2/XA5/MN1/a_324_n18# 0 0.15fF
C7712 XA2/XA5/MP3/a_216_n18# 0 0.03fF
C7713 XA2/CN0 0 3.11fF
C7714 XA2/XA5/MP2/a_216_n18# 0 0.02fF
C7715 XA2/XA5/MP1/a_216_n18# 0 0.03fF
C7716 XA2/XA4/A 0 1.93fF
C7717 XA2/XA4/MN3/a_324_n18# 0 0.15fF
C7718 XA2/XA5/MN0/a_324_n18# 0 0.17fF
C7719 XA2/XA4/MN2/a_324_n18# 0 0.15fF
C7720 XA2/XA4/MN1/a_324_n18# 0 0.15fF
C7721 XA2/XA4/MP3/a_216_n18# 0 0.03fF
C7722 XA2/XA5/MP0/a_216_n18# 0 0.05fF
C7723 XA2/XA4/MP2/a_216_n18# 0 0.02fF
C7724 XA2/XA4/MP1/a_216_n18# 0 0.03fF
C7725 XA2/CN1 0 4.56fF
C7726 XA2/XA3/MN3/a_324_n18# 0 0.15fF
C7727 XA2/XA4/MN0/a_324_n18# 0 0.17fF
C7728 XA2/XA3/MN2/a_324_n18# 0 0.15fF
C7729 XA2/XA3/MN1/a_324_n18# 0 0.15fF
C7730 XA2/XA3/MP3/a_216_n18# 0 0.03fF
C7731 XA2/XA4/MP0/a_216_n18# 0 0.05fF
C7732 D<6> 0 3.91fF
C7733 XA2/XA3/MN0/a_324_n18# 0 0.17fF
C7734 XA2/XA3/MP2/a_216_n18# 0 0.02fF
C7735 XA2/XA3/MP1/a_216_n18# 0 0.03fF
C7736 XA2/XA3/MP0/a_216_n18# 0 0.05fF
C7737 XA2/XA2/A 0 1.31fF
C7738 XA2/XA2/MN3/a_324_n18# 0 0.15fF
C7739 XA2/XA2/MN2/a_324_n18# 0 0.15fF
C7740 XA2/XA2/MN1/a_324_n18# 0 0.15fF
C7741 XA2/XA2/MP3/a_216_n18# 0 0.03fF
C7742 XA2/XA2/MP2/a_216_n18# 0 0.02fF
C7743 XA2/XA2/MP1/a_216_n18# 0 0.03fF
C7744 XA2/XA1/XA5/MN2/S 0 0.06fF
C7745 XA2/XA2/MN0/a_324_n18# 0 0.17fF
C7746 XA2/XA1/XA5/MN1/S 0 0.06fF
C7747 XA2/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7748 XA2/XA1/XA5/MP2/S 0 0.02fF
C7749 XA2/XA2/MP0/a_216_n18# 0 0.05fF
C7750 XA2/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7751 XA2/XA1/XA5/MP1/S 0 0.02fF
C7752 XA2/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7753 XA2/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7754 XA2/XA1/XA4/MN2/S 0 0.06fF
C7755 XA2/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7756 XA2/XA1/XA4/MN1/S 0 0.06fF
C7757 XA2/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7758 XA2/XA1/XA4/MP2/S 0 0.02fF
C7759 XA2/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7760 XA2/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7761 XA2/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7762 XA2/XA1/XA4/MP1/S 0 0.02fF
C7763 XA2/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7764 XA2/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7765 XA2/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7766 XA2/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7767 XA2/XA1/XA2/Y 0 0.78fF
C7768 XA2/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7769 XA2/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7770 XA2/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7771 XA2/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7772 XA2/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7773 XA2/XA1/XA1/MP3/G 0 0.62fF
C7774 XA2/XA1/XA1/MN2/S 0 0.16fF
C7775 XA2/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7776 XA2/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7777 XA3/EN 0 2.02fF
C7778 XA2/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7779 XA2/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7780 XA2/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7781 XA2/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7782 XA2/XA13/MN1/a_324_n18# 0 0.17fF
C7783 XA2/XA13/MN1/a_324_334# 0 0.32fF
C7784 XA2/XA13/MP1/a_216_n18# 0 0.03fF
C7785 XA2/XA13/MP1/a_216_334# 0 0.21fF
C7786 XA2/XA12/MN0/a_324_n18# 0 0.17fF
C7787 XA2/CEO 0 0.35fF
C7788 XA2/XA12/MP0/a_216_n18# 0 0.03fF
C7789 XA2/XA11/MN1/a_324_n18# 0 0.15fF
C7790 XA2/XA11/MP1/S 0 0.02fF
C7791 XA2/XA12/A 0 0.51fF
C7792 XA2/XA11/A 0 0.45fF
C7793 XA2/XA11/MP1/a_216_n18# 0 0.04fF
C7794 XA2/XA9/MN1/a_324_334# 0 0.17fF
C7795 XA2/XA11/MN0/a_324_n18# 0 0.17fF
C7796 XA2/XA9/MP1/a_216_334# 0 0.03fF
C7797 XA2/XA11/MP0/a_216_n18# 0 0.03fF
C7798 XA1/XA9/MN1/S 0 0.05fF
C7799 XA1/XA9/MN1/a_324_n18# 0 0.15fF
C7800 XA1/XA9/Y 0 0.48fF
C7801 XA1/XA9/A 0 0.74fF
C7802 XA1/XA9/MP1/a_216_n18# 0 0.04fF
C7803 XA1/XA9/MN0/a_324_n18# 0 0.17fF
C7804 XA1/DONE 0 0.07fF
C7805 XA1/XA9/MP0/a_216_n18# 0 0.03fF
C7806 XA1/XA7/MN0/a_324_n18# 0 0.17fF
C7807 XA1/XA8/MN0/a_324_n18# 0 0.17fF
C7808 XA1/XA7/MP0/a_216_n18# 0 0.03fF
C7809 XA1/XA8/MP0/a_216_n18# 0 0.02fF
C7810 XA1/XA6/MN3/a_324_n18# 0 0.15fF
C7811 XA1/XA6/MN3/S 0 0.04fF
C7812 XA1/XA6/MN2/a_324_n18# 0 0.15fF
C7813 XA1/XA6/MN1/a_324_n18# 0 0.15fF
C7814 XA1/XA6/MP3/a_216_n18# 0 0.03fF
C7815 XA1/XA6/MN1/S 0 0.04fF
C7816 XA1/XA6/MN0/a_324_n18# 0 0.17fF
C7817 XA1/XA6/MP3/S 0 0.01fF
C7818 XA1/XA6/MP2/a_216_n18# 0 0.02fF
C7819 XA1/XA6/MP1/a_216_n18# 0 0.03fF
C7820 XA1/XA9/B 0 0.83fF
C7821 XA1/XA6/MP1/S 0 0.01fF
C7822 XA1/XA6/MP0/a_216_n18# 0 0.05fF
C7823 XA1/XA5/MN3/a_324_n18# 0 0.15fF
C7824 XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7825 XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7826 XA1/XA5/MP3/a_216_n18# 0 0.03fF
C7827 XA1/XA5/MP2/a_216_n18# 0 0.02fF
C7828 XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7829 XA1/XA4/A 0 1.93fF
C7830 XA1/XA4/MN3/a_324_n18# 0 0.15fF
C7831 XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7832 XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7833 XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7834 XA1/XA4/MP3/a_216_n18# 0 0.03fF
C7835 XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7836 XA1/XA4/MP2/a_216_n18# 0 0.02fF
C7837 XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7838 XA1/XA3/MN3/a_324_n18# 0 0.15fF
C7839 XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7840 XA1/XA3/MN2/a_324_n18# 0 0.15fF
C7841 XA1/XA3/MN1/a_324_n18# 0 0.15fF
C7842 XA1/XA3/MP3/a_216_n18# 0 0.03fF
C7843 XA1/XA4/MP0/a_216_n18# 0 0.05fF
C7844 XA1/XA3/MN0/a_324_n18# 0 0.17fF
C7845 XA1/XA3/MP2/a_216_n18# 0 0.02fF
C7846 XA1/XA3/MP1/a_216_n18# 0 0.03fF
C7847 XA1/XA3/MP0/a_216_n18# 0 0.05fF
C7848 XA1/XA2/A 0 1.31fF
C7849 XA1/XA2/MN3/a_324_n18# 0 0.15fF
C7850 XA1/XA2/MN2/a_324_n18# 0 0.15fF
C7851 XA1/XA2/MN1/a_324_n18# 0 0.15fF
C7852 XA1/XA2/MP3/a_216_n18# 0 0.03fF
C7853 XA1/XA2/MP2/a_216_n18# 0 0.02fF
C7854 XA1/XA2/MP1/a_216_n18# 0 0.03fF
C7855 XA1/XA1/XA5/MN2/S 0 0.06fF
C7856 XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7857 XA1/XA1/XA5/MN1/S 0 0.06fF
C7858 XA1/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C7859 XA1/XA1/XA5/MP2/S 0 0.02fF
C7860 XA1/XA2/MP0/a_216_n18# 0 0.05fF
C7861 XA1/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C7862 XA1/XA1/XA5/MP1/S 0 0.02fF
C7863 XA1/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C7864 XA1/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C7865 XA1/XA1/XA4/MN2/S 0 0.06fF
C7866 XA1/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C7867 XA1/XA1/XA4/MN1/S 0 0.06fF
C7868 XA1/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C7869 XA1/XA1/XA4/MP2/S 0 0.02fF
C7870 XA1/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C7871 XA1/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C7872 XA1/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C7873 XA1/XA1/XA4/MP1/S 0 0.02fF
C7874 XA1/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C7875 XA1/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C7876 XA1/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C7877 XA1/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C7878 XA1/XA1/XA2/Y 0 0.78fF
C7879 XA1/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C7880 XA1/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C7881 XA1/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C7882 XA1/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C7883 XA1/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C7884 XA1/XA1/XA1/MP3/G 0 0.62fF
C7885 XA1/XA1/XA1/MN2/S 0 0.16fF
C7886 XA1/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C7887 XA1/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C7888 XA2/EN 0 2.13fF
C7889 XA1/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C7890 XA1/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C7891 XA1/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C7892 XA1/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C7893 XA1/XA13/MN1/a_324_n18# 0 0.17fF
C7894 XA1/XA13/MN1/a_324_334# 0 0.32fF
C7895 XA1/XA13/MP1/a_216_n18# 0 0.03fF
C7896 XA1/XA13/MP1/a_216_334# 0 0.21fF
C7897 XA1/XA12/MN0/a_324_n18# 0 0.17fF
C7898 XA1/CEO 0 0.58fF
C7899 XA1/XA12/MP0/a_216_n18# 0 0.03fF
C7900 XA1/XA11/MN1/a_324_n18# 0 0.15fF
C7901 XA1/XA11/MP1/S 0 0.02fF
C7902 XA1/XA12/A 0 0.51fF
C7903 XA1/XA11/A 0 0.45fF
C7904 XA1/XA11/MP1/a_216_n18# 0 0.04fF
C7905 XA1/XA9/MN1/a_324_334# 0 0.17fF
C7906 XA1/XA11/MN0/a_324_n18# 0 0.17fF
C7907 XA1/XA9/MP1/a_216_334# 0 0.03fF
C7908 XA1/XA11/MP0/a_216_n18# 0 0.03fF
C7909 XB2/XA7/MN1/a_324_n18# 0 0.17fF
C7910 XB2/XA7/MP1/a_216_n18# 0 0.02fF
C7911 XB2/XA5b/MN1/a_324_n18# 0 0.32fF
C7912 XB2/XA0/MN0/a_324_n18# 0 0.17fF
C7913 XB2/XA5b/MP1/a_216_n18# 0 0.21fF
C7914 XB2/XA0/MP0/a_216_n18# 0 0.03fF
C7915 XB2/XA4/MN1/S 0 0.05fF
C7916 XB2/XA1/Y 0 0.35fF
C7917 XB2/XA4/MN1/a_324_334# 0 0.17fF
C7918 XB2/XA4/MN0/a_324_n18# 0 0.17fF
C7919 XB2/XA4/MN1/a_324_n18# 0 0.15fF
C7920 XB2/XA4/GNG 0 67.61fF
C7921 XB2/XA4/MP1/a_216_334# 0 0.03fF
C7922 XB2/XA4/MP0/a_216_n18# 0 0.04fF
C7923 XB2/XA4/MP1/a_216_n18# 0 0.04fF
C7924 XB2/XA5/MN1/a_324_334# 0 0.32fF
C7925 XB2/XA5/MP1/a_216_334# 0 0.21fF
C7926 XB2/XA3/MN2/a_324_n18# 0 0.15fF
C7927 XB2/XA3/B 0 71.43fF
C7928 XB2/XA3/MN1/a_324_n18# 0 0.15fF
C7929 XB2/XA3/MP0/S 0 0.64fF
C7930 XB2/XA3/MN0/a_324_n18# 0 0.17fF
C7931 XB2/XA3/MP2/a_216_n18# 0 0.03fF
C7932 XB2/XA3/MP0/a_216_n18# 0 0.04fF
C7933 XB2/XA3/MP0/a_216_334# 0 0.03fF
C7934 XB2/XA7/MN1/a_324_334# 0 0.17fF
C7935 XB2/XA5/MN1/a_324_n18# 0 0.17fF
C7936 XB2/XA2/MP0/G 0 0.52fF
C7937 XB2/XA7/MP1/a_216_334# 0 0.03fF
C7938 XB2/XA5/MP1/a_216_n18# 0 0.03fF
C7939 XB2/XA1/MP0/G 0 0.56fF
C7940 XB2/CKN 0 1.12fF
C7941 XB2/M8/a_324_n18# 0 0.16fF
C7942 XB2/M8/a_324_334# 0 0.32fF
C7943 XB2/M7/a_324_n18# 0 0.16fF
C7944 XB2/M6/a_324_n18# 0 0.16fF
C7945 XB2/M5/a_324_n18# 0 0.16fF
C7946 XB2/M3/a_324_n18# 0 0.16fF
C7947 XB2/M4/a_324_n18# 0 0.16fF
C7948 XB2/M2/a_324_n18# 0 0.16fF
C7949 SAR_IN 0 1.04fF
C7950 XB2/M4/G 0 1.49fF
C7951 XB2/M1/a_324_n18# 0 0.32fF
C7952 XA0/XA9/MN1/S 0 0.05fF
C7953 XA0/XA9/MN1/a_324_n18# 0 0.15fF
C7954 XA0/XA9/Y 0 0.48fF
C7955 XA0/XA9/A 0 0.74fF
C7956 XA0/XA9/MP1/a_216_n18# 0 0.04fF
C7957 XA0/XA9/MN0/a_324_n18# 0 0.17fF
C7958 XA0/DONE 0 0.07fF
C7959 XA0/XA9/MP0/a_216_n18# 0 0.03fF
C7960 XA0/XA7/MN0/a_324_n18# 0 0.17fF
C7961 XA0/XA8/MN0/a_324_n18# 0 0.17fF
C7962 XA0/XA7/MP0/a_216_n18# 0 0.03fF
C7963 XA0/XA8/MP0/a_216_n18# 0 0.02fF
C7964 XA0/XA6/MN3/a_324_n18# 0 0.15fF
C7965 XA0/XA6/MN3/S 0 0.04fF
C7966 XA0/XA6/MN2/a_324_n18# 0 0.15fF
C7967 XA0/XA6/MN1/a_324_n18# 0 0.15fF
C7968 XA0/XA6/MP3/a_216_n18# 0 0.03fF
C7969 CK_SAMPLE 0 8.64fF
C7970 XA0/XA6/MN1/S 0 0.04fF
C7971 XA0/XA6/MN0/a_324_n18# 0 0.17fF
C7972 XA0/XA6/MP3/S 0 0.01fF
C7973 XA0/XA6/MP2/a_216_n18# 0 0.02fF
C7974 XA0/XA6/MP1/a_216_n18# 0 0.03fF
C7975 XA0/XA9/B 0 0.83fF
C7976 XA0/XA6/MP1/S 0 0.01fF
C7977 XA0/XA6/MP0/a_216_n18# 0 0.05fF
C7978 XA0/XA5/MN3/a_324_n18# 0 0.15fF
C7979 XA0/XA5/MN2/a_324_n18# 0 0.15fF
C7980 XA0/XA5/MN1/a_324_n18# 0 0.15fF
C7981 XA0/XA5/MP3/a_216_n18# 0 0.03fF
C7982 XA0/XA5/MP2/a_216_n18# 0 0.02fF
C7983 XA0/XA5/MP1/a_216_n18# 0 0.03fF
C7984 XA0/XA4/A 0 1.93fF
C7985 XA0/XA4/MN3/a_324_n18# 0 0.15fF
C7986 XA0/XA5/MN0/a_324_n18# 0 0.17fF
C7987 XA0/XA4/MN2/a_324_n18# 0 0.15fF
C7988 XA0/XA4/MN1/a_324_n18# 0 0.15fF
C7989 XA0/XA4/MP3/a_216_n18# 0 0.03fF
C7990 XA0/XA5/MP0/a_216_n18# 0 0.05fF
C7991 XA0/XA4/MP2/a_216_n18# 0 0.02fF
C7992 XA0/XA4/MP1/a_216_n18# 0 0.03fF
C7993 XA0/XA3/MN3/a_324_n18# 0 0.15fF
C7994 XA0/XA4/MN0/a_324_n18# 0 0.17fF
C7995 XA0/XA3/MN2/a_324_n18# 0 0.15fF
C7996 XA0/XA3/MN1/a_324_n18# 0 0.15fF
C7997 XA0/XA3/MP3/a_216_n18# 0 0.03fF
C7998 XA0/XA4/MP0/a_216_n18# 0 0.05fF
C7999 XA0/XA3/MN0/a_324_n18# 0 0.17fF
C8000 XA0/XA3/MP2/a_216_n18# 0 0.02fF
C8001 XA0/XA3/MP1/a_216_n18# 0 0.03fF
C8002 XA0/XA3/MP0/a_216_n18# 0 0.05fF
C8003 XA0/XA2/A 0 1.31fF
C8004 XA0/XA2/MN3/a_324_n18# 0 0.15fF
C8005 XA0/XA2/MN2/a_324_n18# 0 0.15fF
C8006 XA0/XA2/MN1/a_324_n18# 0 0.15fF
C8007 XA0/XA2/MP3/a_216_n18# 0 0.03fF
C8008 XA0/XA2/MP2/a_216_n18# 0 0.02fF
C8009 VREF 0 33.40fF
C8010 XA0/XA2/MP1/a_216_n18# 0 0.03fF
C8011 EN 0 3.06fF
C8012 XA0/XA1/XA5/MN2/S 0 0.06fF
C8013 XA0/XA2/MN0/a_324_n18# 0 0.17fF
C8014 XA0/XA1/XA5/MN1/S 0 0.06fF
C8015 XA0/XA1/XA5/MN2/a_324_n18# 0 0.15fF
C8016 XA0/XA1/XA5/MP2/S 0 0.02fF
C8017 XA0/XA2/MP0/a_216_n18# 0 0.05fF
C8018 XA0/XA1/XA5/MN1/a_324_n18# 0 0.15fF
C8019 XA0/XA1/XA5/MP1/S 0 0.02fF
C8020 XA0/XA1/XA5/MP2/a_216_n18# 0 0.03fF
C8021 XA0/XA1/XA5/MP1/a_216_n18# 0 0.03fF
C8022 XA0/XA1/XA4/MN2/S 0 0.06fF
C8023 XA0/XA1/XA5/MN0/a_324_n18# 0 0.17fF
C8024 XA0/XA1/XA4/MN1/S 0 0.06fF
C8025 XA0/XA1/XA4/MN2/a_324_n18# 0 0.15fF
C8026 XA0/XA1/XA4/MP2/S 0 0.02fF
C8027 XA0/XA1/XA5/MP0/a_216_n18# 0 0.05fF
C8028 XA0/XA1/XA4/MN0/a_324_n18# 0 0.17fF
C8029 XA0/XA1/XA4/MN1/a_324_n18# 0 0.15fF
C8030 XA0/XA1/XA4/MP1/S 0 0.02fF
C8031 XA0/XA1/XA4/MP2/a_216_n18# 0 0.03fF
C8032 XA0/XA1/XA4/MP0/a_216_n18# 0 0.03fF
C8033 XA0/XA1/XA4/MP1/a_216_n18# 0 0.03fF
C8034 XA0/XA1/XA2/MN0/a_324_n18# 0 0.17fF
C8035 XA0/XA1/XA2/Y 0 0.78fF
C8036 XA0/XA1/XA2/MP0/a_216_n18# 0 0.03fF
C8037 XA20/CNO 0 8.06fF
C8038 XA20/CPO 0 6.87fF
C8039 XA0/XA1/XA1/MN3/a_324_n18# 0 0.15fF
C8040 XA0/XA1/XA1/MN2/a_324_n18# 0 0.15fF
C8041 XA0/XA1/XA1/MN1/a_324_n18# 0 0.15fF
C8042 XA0/XA1/XA1/MP3/a_216_n18# 0 0.03fF
C8043 XA0/XA1/XA1/MP3/G 0 0.62fF
C8044 XA0/XA1/XA1/MN2/S 0 0.16fF
C8045 XA0/XA1/XA1/MN0/a_324_n18# 0 0.17fF
C8046 XA0/XA1/XA1/MP2/a_216_n18# 0 0.02fF
C8047 XA1/EN 0 2.19fF
C8048 XA0/XA1/XA1/MP1/a_216_n18# 0 0.03fF
C8049 XA0/XA1/XA1/MP0/a_216_n18# 0 0.05fF
C8050 XA0/XA1/XA0/MN1/a_324_n18# 0 0.32fF
C8051 AVDD 0 747.75fF
C8052 XA0/XA1/XA0/MP1/a_216_n18# 0 0.21fF
C8053 XA0/XA13/MN1/a_324_n18# 0 0.17fF
C8054 XA0/XA13/MN1/a_324_334# 0 0.32fF
C8055 XA0/XA13/MP1/a_216_n18# 0 0.03fF
C8056 XA0/XA13/MP1/a_216_334# 0 0.21fF
C8057 XA0/XA12/MN0/a_324_n18# 0 0.17fF
C8058 XA0/CEO 0 0.39fF
C8059 XA0/XA12/MP0/a_216_n18# 0 0.03fF
C8060 XA0/XA11/MN1/a_324_n18# 0 0.15fF
C8061 XA0/XA11/MP1/S 0 0.02fF
C8062 XA0/XA12/A 0 0.51fF
C8063 XA0/XA11/A 0 0.45fF
C8064 XA0/XA11/MP1/a_216_n18# 0 0.04fF
C8065 XA0/XA9/MN1/a_324_334# 0 0.17fF
C8066 XA0/XA11/MN0/a_324_n18# 0 0.17fF
C8067 XA0/XA9/MP1/a_216_334# 0 0.03fF
C8068 XA0/XA11/MP0/a_216_n18# 0 0.03fF
C8069 XB1/XA7/MN1/a_324_n18# 0 0.17fF
C8070 XB1/XA7/MP1/a_216_n18# 0 0.02fF
C8071 AVSS 0 258.84fF
C8072 XB1/XA5b/MN1/a_324_n18# 0 0.32fF
C8073 XB1/XA0/MN0/a_324_n18# 0 0.17fF
C8074 XB1/XA5b/MP1/a_216_n18# 0 0.21fF
C8075 XB1/XA0/MP0/a_216_n18# 0 0.03fF
C8076 XB1/XA4/MN1/S 0 0.05fF
C8077 XB1/XA1/Y 0 0.35fF
C8078 XB1/XA4/MN1/a_324_334# 0 0.17fF
C8079 XB1/XA4/MN0/a_324_n18# 0 0.17fF
C8080 XB1/XA4/MN1/a_324_n18# 0 0.15fF
C8081 XB1/XA4/GNG 0 67.61fF
C8082 XB1/XA4/MP1/a_216_334# 0 0.03fF
C8083 XB1/XA4/MP0/a_216_n18# 0 0.04fF
C8084 XB1/XA4/MP1/a_216_n18# 0 0.04fF
C8085 XB1/XA5/MN1/a_324_334# 0 0.32fF
C8086 XB1/XA5/MP1/a_216_334# 0 0.21fF
C8087 XB1/XA3/MN2/a_324_n18# 0 0.15fF
C8088 XB1/XA3/B 0 71.43fF
C8089 XB1/XA3/MN1/a_324_n18# 0 0.15fF
C8090 XB1/XA3/MP0/S 0 0.64fF
C8091 XB1/XA3/MN0/a_324_n18# 0 0.17fF
C8092 XB1/XA3/MP2/a_216_n18# 0 0.03fF
C8093 XB1/XA3/MP0/a_216_n18# 0 0.04fF
C8094 XB1/XA3/MP0/a_216_334# 0 0.03fF
C8095 XB1/XA7/MN1/a_324_334# 0 0.17fF
C8096 XB1/XA5/MN1/a_324_n18# 0 0.17fF
C8097 XB1/XA2/MP0/G 0 0.52fF
C8098 XB1/XA7/MP1/a_216_334# 0 0.03fF
C8099 XB1/XA5/MP1/a_216_n18# 0 0.03fF
C8100 XB1/XA1/MP0/G 0 0.56fF
C8101 CK_SAMPLE_BSSW 0 2.77fF
C8102 XB1/CKN 0 1.12fF
C8103 XB1/M8/a_324_n18# 0 0.16fF
C8104 XB1/M8/a_324_334# 0 0.32fF
C8105 XB1/M7/a_324_n18# 0 0.16fF
C8106 XB1/M6/a_324_n18# 0 0.16fF
C8107 XA0/CEIN 0 21.38fF
C8108 XB1/M5/a_324_n18# 0 0.16fF
C8109 XB1/M3/a_324_n18# 0 0.16fF
C8110 XB1/M4/a_324_n18# 0 0.16fF
C8111 XB1/M2/a_324_n18# 0 0.16fF
C8112 SAR_IP 0 0.99fF
C8113 XB1/M4/G 0 1.49fF
C8114 SARP 0 17.29fF
C8115 XB1/M1/a_324_n18# 0 0.32fF
C8116 XA20/XA9/MN0/a_324_n18# 0 0.17fF
C8117 XA20/XA9/MP0/a_216_n18# 0 0.03fF
C8118 XA20/XA3/CO 0 1.52fF
C8119 XA20/XA2a/MN3/a_324_n18# 0 0.15fF
C8120 XA20/XA2a/MN2/a_324_n18# 0 0.15fF
C8121 XA20/XA2a/MN1/a_324_n18# 0 0.15fF
C8122 XA20/XA2a/MP3/a_216_n18# 0 0.03fF
C8123 XA20/XA2/MN6/a_324_334# 0 0.17fF
C8124 XA20/XA2a/MP2/a_216_n18# 0 0.02fF
C8125 XA20/XA2a/MP1/a_216_n18# 0 0.03fF
C8126 XA20/XA2/MP6/a_216_334# 0 0.05fF
C8127 XA20/XA3a/A 0 1.71fF
C8128 XA20/XA3a/MN3/a_324_n18# 0 0.15fF
C8129 XA20/XA3/MN0/a_324_n18# 0 0.17fF
C8130 XA20/XA3a/MN2/a_324_n18# 0 0.15fF
C8131 XA20/XA3a/MN1/a_324_n18# 0 0.15fF
C8132 XA20/XA3a/MP3/a_216_n18# 0 0.03fF
C8133 XA20/XA3/MP0/a_216_n18# 0 0.05fF
C8134 XA20/XA3a/MN0/a_324_n18# 0 0.17fF
C8135 XA20/XA3a/MP2/a_216_n18# 0 0.02fF
C8136 XA20/XA3a/MP1/a_216_n18# 0 0.03fF
C8137 XA20/XA3a/MP0/a_216_n18# 0 0.05fF
C8138 XA20/XA4/MP5_DMY/a_216_n18# 0 0.02fF
C8139 XA20/XA4/MP2_DMY/a_216_n18# 0 0.02fF
C8140 XA20/XA4/MP6_DMY/a_216_n18# 0 0.02fF
C8141 XA20/XA4/MP3_DMY/a_216_n18# 0 0.01fF
C8142 XA20/XA4/MN5/a_324_n18# 0 0.15fF
C8143 XA20/XA4/MN6/a_324_n18# 0 0.15fF
C8144 XA20/XA4/MN4/a_324_n18# 0 0.15fF
C8145 XA20/XA4/MN3/a_324_n18# 0 0.15fF
C8146 XA20/XA4/MN2/a_324_n18# 0 0.15fF
C8147 XA20/XA4/MN1/a_324_n18# 0 0.15fF
C8148 XA20/XA4/MP0/S 0 0.47fF
C8149 XA20/XA4/MN0/a_324_n18# 0 0.17fF
C8150 XA20/XA4/MP0/a_216_n18# 0 0.05fF
C8151 XA20/XA4/MP4_DMY/a_216_n18# 0 0.01fF
C8152 XA20/XA4/MP0/a_216_334# 0 0.02fF
C8153 XA20/XA3/MN5/a_324_n18# 0 0.15fF
C8154 XA20/XA3/MN6/a_324_n18# 0 0.15fF
C8155 XA20/XA3/MN4/a_324_n18# 0 0.15fF
C8156 XA20/XA3/MP6/a_216_n18# 0 0.02fF
C8157 XA20/XA3/MN3/a_324_n18# 0 0.15fF
C8158 XA20/XA3/MP5/a_216_n18# 0 0.02fF
C8159 XA20/XA3/MN2/a_324_n18# 0 0.15fF
C8160 XA20/XA3/MP4/a_216_n18# 0 0.01fF
C8161 XA20/XA3/N2 0 0.35fF
C8162 XA20/XA3/MN1/a_324_n18# 0 0.15fF
C8163 XA20/XA3/MP3/a_216_n18# 0 0.01fF
C8164 XA20/XA3/MP2/a_216_n18# 0 0.02fF
C8165 XA20/XA3/MP1/a_216_n18# 0 0.02fF
C8166 XA20/XA9/Y 0 2.27fF
C8167 XA20/XA2/MN5/a_324_n18# 0 0.15fF
C8168 XA20/XA2/MN6/a_324_n18# 0 0.15fF
C8169 XA20/XA2/MN4/a_324_n18# 0 0.15fF
C8170 XA20/XA2/MP6/a_216_n18# 0 0.02fF
C8171 XA20/XA2/MN3/a_324_n18# 0 0.15fF
C8172 XA20/XA2/MP5/a_216_n18# 0 0.02fF
C8173 XA20/XA2/MN2/a_324_n18# 0 0.15fF
C8174 XA20/XA2/MP4/a_216_n18# 0 0.01fF
C8175 XA20/XA2/N2 0 0.35fF
C8176 XA20/XA2/MN1/a_324_n18# 0 0.15fF
C8177 XA20/XA2/MP3/a_216_n18# 0 0.01fF
C8178 XA20/XA3/N1 0 0.97fF
C8179 XA20/XA2/MN0/a_324_n18# 0 0.17fF
C8180 XA20/XA2/MP2/a_216_n18# 0 0.02fF
C8181 XA20/XA2/MP1/a_216_n18# 0 0.02fF
C8182 XA20/XA2/MP0/a_216_n18# 0 0.05fF
C8183 XA20/XA9/A 0 2.65fF
C8184 XA20/XA1/MP5_DMY/a_216_n18# 0 0.02fF
C8185 XA20/XA1/MP2_DMY/a_216_n18# 0 0.02fF
C8186 XA20/XA1/MP6_DMY/a_216_n18# 0 0.02fF
C8187 XA20/XA1/MP3_DMY/a_216_n18# 0 0.01fF
C8188 XA20/XA1/MN5/a_324_n18# 0 0.15fF
C8189 XA20/XA1/MN6/a_324_n18# 0 0.15fF
C8190 XA20/XA1/MN4/a_324_n18# 0 0.15fF
C8191 XA20/XA1/MN3/a_324_n18# 0 0.15fF
C8192 XA20/XA1/MN2/a_324_n18# 0 0.15fF
C8193 XA20/XA1/MN1/a_324_n18# 0 0.15fF
C8194 XA20/XA1/MP0/S 0 0.47fF
C8195 XA20/XA1/MN0/a_324_n18# 0 0.17fF
C8196 XA20/XA1/MP0/a_216_n18# 0 0.05fF
C8197 XA20/XA1/MP4_DMY/a_216_n18# 0 0.01fF
C8198 XA20/XA1/MP0/a_216_334# 0 0.02fF
C8199 XA20/XA0/MN1/a_324_n18# 0 0.32fF
C8200 XA20/XA0/MP1/a_216_n18# 0 0.21fF
C8201 XA20/XA13/MN1/a_324_334# 0 0.32fF
C8202 XA20/XA13/MP1/a_216_334# 0 0.21fF
C8203 XA20/XA13/MN1/a_324_n18# 0 0.17fF
C8204 XA20/XA13/MP1/a_216_n18# 0 0.03fF
C8205 XA20/XA12/MN0/a_324_n18# 0 0.17fF
C8206 XA20/XA11/MN0/a_324_n18# 0 0.17fF
C8207 XA20/XA11/MN1/a_324_n18# 0 0.15fF
C8208 XA20/XA11/MP1/S 0 0.02fF
C8209 XA20/XA12/MP0/a_216_n18# 0 0.03fF
C8210 XA20/XA11/MP0/a_216_n18# 0 0.03fF
C8211 XA20/XA11/MP1/a_216_n18# 0 0.04fF
C8212 XA20/XA10/MN1/S 0 0.05fF
C8213 XA20/XA9/MN0/a_324_334# 0 0.17fF
C8214 XA20/XA10/MN1/a_324_n18# 0 0.15fF
C8215 XA20/XA12/Y 0 0.38fF
C8216 XA20/XA11/Y 0 0.58fF
C8217 XA20/XA9/MP0/a_216_334# 0 0.03fF
C8218 XA20/XA10/MP1/a_216_n18# 0 0.04fF
C8219 XA0/CN0 0 8.47fF
C8220 XA1/CN0 0 4.41fF
C8221 D<8> 0 7.01fF
C8222 XA3/CN1 0 4.39fF
C8223 XA1/CN1 0 4.45fF
C8224 XDAC2/XC32a<0>/XRES16/B 0 2.89fF
C8225 XDAC2/XC32a<0>/XRES8/B 0 1.96fF
C8226 XDAC2/XC32a<0>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8227 XDAC2/XC32a<0>/XRES4/B 0 1.62fF
C8228 XDAC2/XC32a<0>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8229 XDAC2/XC32a<0>/XRES1B/B 0 2.43fF
C8230 XDAC2/XC32a<0>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8231 XDAC2/XC32a<0>/XRES2/B 0 1.42fF
C8232 XDAC2/XC32a<0>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8233 XDAC2/XC32a<0>/C1A 0 0.09fF
C8234 XDAC2/XC32a<0>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8235 XDAC2/XC32a<0>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8236 XDAC2/XC128a<1>/XRES16/B 0 2.89fF
C8237 XDAC2/XC128a<1>/XRES8/B 0 1.96fF
C8238 XDAC2/XC128a<1>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8239 XDAC2/XC128a<1>/XRES4/B 0 1.62fF
C8240 XDAC2/XC128a<1>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8241 XDAC2/XC128a<1>/XRES1B/B 0 2.43fF
C8242 XDAC2/XC128a<1>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8243 XDAC2/XC128a<1>/XRES2/B 0 1.42fF
C8244 XDAC2/XC128a<1>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8245 XDAC2/XC128a<1>/XRES1A/B 0 1.29fF
C8246 XDAC2/XC128a<1>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8247 XDAC2/XC128a<1>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8248 XDAC2/XC64b<1>/XRES16/B 0 2.89fF
C8249 XDAC2/XC64b<1>/XRES8/B 0 1.96fF
C8250 XDAC2/XC64b<1>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8251 XDAC2/XC64b<1>/XRES4/B 0 1.62fF
C8252 XDAC2/XC64b<1>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8253 XDAC2/XC64b<1>/XRES1B/B 0 2.43fF
C8254 XDAC2/XC64b<1>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8255 XDAC2/XC64b<1>/XRES2/B 0 1.42fF
C8256 XDAC2/XC64b<1>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8257 XDAC2/XC64b<1>/XRES1A/B 0 1.29fF
C8258 XDAC2/XC64b<1>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8259 XDAC2/XC64b<1>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8260 XDAC2/XC1/XRES16/B 0 2.89fF
C8261 XDAC2/XC1/XRES8/B 0 1.96fF
C8262 XDAC2/XC1/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8263 XDAC2/XC1/XRES4/B 0 1.62fF
C8264 XDAC2/XC1/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8265 XDAC2/XC1/XRES1B/B 0 2.43fF
C8266 XDAC2/XC1/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8267 XDAC2/XC1/XRES2/B 0 1.42fF
C8268 XDAC2/XC1/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8269 XDAC2/XC1/XRES1A/B 0 1.29fF
C8270 XDAC2/XC1/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8271 XDAC2/XC1/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8272 XDAC2/XC0/XRES16/B 0 2.89fF
C8273 XDAC2/XC0/XRES8/B 0 1.96fF
C8274 XDAC2/XC0/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8275 XDAC2/XC0/XRES4/B 0 1.62fF
C8276 XDAC2/XC0/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8277 XDAC2/XC0/XRES1B/B 0 2.43fF
C8278 XDAC2/XC0/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8279 XDAC2/XC0/XRES2/B 0 1.42fF
C8280 XDAC2/XC0/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8281 XDAC2/XC0/XRES1A/B 0 1.29fF
C8282 XDAC2/XC0/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8283 XDAC2/XC0/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8284 SARN 0 19.23fF
C8285 XDAC2/XC64a<0>/XRES16/B 0 2.89fF
C8286 XDAC2/XC64a<0>/XRES8/B 0 1.96fF
C8287 XDAC2/XC64a<0>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8288 XDAC2/XC64a<0>/XRES4/B 0 1.62fF
C8289 XDAC2/XC64a<0>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8290 XDAC2/XC64a<0>/XRES1B/B 0 2.43fF
C8291 XDAC2/XC64a<0>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8292 XDAC2/XC64a<0>/XRES2/B 0 1.42fF
C8293 XDAC2/XC64a<0>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8294 XDAC2/XC64a<0>/XRES1A/B 0 1.29fF
C8295 XDAC2/XC64a<0>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8296 XDAC2/XC64a<0>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8297 XDAC2/X16ab/XRES16/B 0 2.89fF
C8298 XDAC2/X16ab/XRES8/B 0 1.96fF
C8299 XDAC2/X16ab/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8300 XDAC2/X16ab/XRES4/B 0 1.62fF
C8301 XDAC2/X16ab/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8302 XDAC2/X16ab/XRES1B/B 0 2.43fF
C8303 XDAC2/X16ab/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8304 XDAC2/X16ab/XRES2/B 0 1.42fF
C8305 XDAC2/X16ab/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8306 XDAC2/X16ab/XRES1A/B 0 1.29fF
C8307 XDAC2/X16ab/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8308 XDAC2/X16ab/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8309 XDAC2/XC128b<2>/XRES16/B 0 2.89fF
C8310 XDAC2/XC128b<2>/XRES8/B 0 1.96fF
C8311 XDAC2/XC128b<2>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8312 XDAC2/XC128b<2>/XRES4/B 0 1.62fF
C8313 XDAC2/XC128b<2>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8314 XDAC2/XC128b<2>/XRES1B/B 0 2.43fF
C8315 XDAC2/XC128b<2>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8316 XDAC2/XC128b<2>/XRES2/B 0 1.42fF
C8317 XDAC2/XC128b<2>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8318 XDAC2/XC128b<2>/XRES1A/B 0 1.29fF
C8319 XDAC2/XC128b<2>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8320 XDAC2/XC128b<2>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8321 XA0/CP0 0 8.68fF
C8322 XA1/CP0 0 6.70fF
C8323 XA0/CP1 0 6.32fF
C8324 D<5> 0 3.31fF
C8325 D<7> 0 3.42fF
C8326 XDAC1/XC32a<0>/XRES16/B 0 2.89fF
C8327 XDAC1/XC32a<0>/XRES8/B 0 1.96fF
C8328 XDAC1/XC32a<0>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8329 XDAC1/XC32a<0>/XRES4/B 0 1.62fF
C8330 XDAC1/XC32a<0>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8331 XDAC1/XC32a<0>/XRES1B/B 0 2.43fF
C8332 XDAC1/XC32a<0>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8333 XDAC1/XC32a<0>/XRES2/B 0 1.42fF
C8334 XDAC1/XC32a<0>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8335 XDAC1/XC32a<0>/C1A 0 0.09fF
C8336 XDAC1/XC32a<0>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8337 XDAC1/XC32a<0>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8338 XDAC1/XC128a<1>/XRES16/B 0 2.89fF
C8339 XDAC1/XC128a<1>/XRES8/B 0 1.96fF
C8340 XDAC1/XC128a<1>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8341 XDAC1/XC128a<1>/XRES4/B 0 1.62fF
C8342 XDAC1/XC128a<1>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8343 XDAC1/XC128a<1>/XRES1B/B 0 2.43fF
C8344 XDAC1/XC128a<1>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8345 XDAC1/XC128a<1>/XRES2/B 0 1.42fF
C8346 XDAC1/XC128a<1>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8347 XDAC1/XC128a<1>/XRES1A/B 0 1.29fF
C8348 XDAC1/XC128a<1>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8349 XDAC1/XC128a<1>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8350 XDAC1/XC64b<1>/XRES16/B 0 2.89fF
C8351 XDAC1/XC64b<1>/XRES8/B 0 1.96fF
C8352 XDAC1/XC64b<1>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8353 XDAC1/XC64b<1>/XRES4/B 0 1.62fF
C8354 XDAC1/XC64b<1>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8355 XDAC1/XC64b<1>/XRES1B/B 0 2.43fF
C8356 XDAC1/XC64b<1>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8357 XDAC1/XC64b<1>/XRES2/B 0 1.42fF
C8358 XDAC1/XC64b<1>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8359 XDAC1/XC64b<1>/XRES1A/B 0 1.29fF
C8360 XDAC1/XC64b<1>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8361 XDAC1/XC64b<1>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8362 XDAC1/XC1/XRES16/B 0 2.89fF
C8363 XDAC1/XC1/XRES8/B 0 1.96fF
C8364 XDAC1/XC1/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8365 XDAC1/XC1/XRES4/B 0 1.62fF
C8366 XDAC1/XC1/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8367 XDAC1/XC1/XRES1B/B 0 2.43fF
C8368 XDAC1/XC1/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8369 XDAC1/XC1/XRES2/B 0 1.42fF
C8370 XDAC1/XC1/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8371 XDAC1/XC1/XRES1A/B 0 1.29fF
C8372 XDAC1/XC1/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8373 XDAC1/XC1/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8374 XDAC1/XC0/XRES16/B 0 2.89fF
C8375 XDAC1/XC0/XRES8/B 0 1.96fF
C8376 XDAC1/XC0/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8377 XDAC1/XC0/XRES4/B 0 1.62fF
C8378 XDAC1/XC0/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8379 XDAC1/XC0/XRES1B/B 0 2.43fF
C8380 XDAC1/XC0/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8381 XDAC1/XC0/XRES2/B 0 1.42fF
C8382 XDAC1/XC0/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8383 XDAC1/XC0/XRES1A/B 0 1.29fF
C8384 XDAC1/XC0/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8385 XDAC1/XC0/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8386 XDAC1/XC64a<0>/XRES16/B 0 2.89fF
C8387 XDAC1/XC64a<0>/XRES8/B 0 1.96fF
C8388 XDAC1/XC64a<0>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8389 XDAC1/XC64a<0>/XRES4/B 0 1.62fF
C8390 XDAC1/XC64a<0>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8391 XDAC1/XC64a<0>/XRES1B/B 0 2.43fF
C8392 XDAC1/XC64a<0>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8393 XDAC1/XC64a<0>/XRES2/B 0 1.42fF
C8394 XDAC1/XC64a<0>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8395 XDAC1/XC64a<0>/XRES1A/B 0 1.29fF
C8396 XDAC1/XC64a<0>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8397 XDAC1/XC64a<0>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8398 XDAC1/X16ab/XRES16/B 0 2.89fF
C8399 XDAC1/X16ab/XRES8/B 0 1.96fF
C8400 XDAC1/X16ab/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8401 XDAC1/X16ab/XRES4/B 0 1.62fF
C8402 XDAC1/X16ab/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8403 XDAC1/X16ab/XRES1B/B 0 2.43fF
C8404 XDAC1/X16ab/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8405 XDAC1/X16ab/XRES2/B 0 1.42fF
C8406 XDAC1/X16ab/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8407 XDAC1/X16ab/XRES1A/B 0 1.29fF
C8408 XDAC1/X16ab/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8409 XDAC1/X16ab/XRES16/li_60_0# 0 0.03fF $ **FLOATING
C8410 XDAC1/XC128b<2>/XRES16/B 0 2.89fF
C8411 XDAC1/XC128b<2>/XRES8/B 0 1.96fF
C8412 XDAC1/XC128b<2>/XRES8/li_60_0# 0 0.03fF $ **FLOATING
C8413 XDAC1/XC128b<2>/XRES4/B 0 1.62fF
C8414 XDAC1/XC128b<2>/XRES4/li_60_0# 0 0.03fF $ **FLOATING
C8415 XDAC1/XC128b<2>/XRES1B/B 0 2.43fF
C8416 XDAC1/XC128b<2>/XRES1B/li_60_0# 0 0.03fF $ **FLOATING
C8417 XDAC1/XC128b<2>/XRES2/B 0 1.42fF
C8418 XDAC1/XC128b<2>/XRES2/li_60_0# 0 0.03fF $ **FLOATING
C8419 XDAC1/XC128b<2>/XRES1A/B 0 1.29fF
C8420 XDAC1/XC128b<2>/XRES1A/li_60_0# 0 0.03fF $ **FLOATING
C8421 XDAC1/XC128b<2>/XRES16/li_60_0# 0 0.03fF $ **FLOATING
.ends
