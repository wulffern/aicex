magic
tech sky130A
magscale 1 2
timestamp 1660667839
<< checkpaint >>
rect -1104 -1104 38440 27024
<< locali >>
rect 38200 -1104 38440 27024
rect -1104 -1104 38440 -864
rect -1104 26784 38440 27024
rect -1104 -1104 -864 27024
rect 38200 -1104 38440 27024
rect -864 -200 -640 -88
rect -864 4380 -640 4492
rect -864 8960 -640 9072
rect -864 13540 -640 13652
rect -864 18120 -640 18232
rect 2106 21510 2430 21730
rect -54 3190 270 3410
<< m3 >>
rect 20348 -1104 20564 40
rect 20456 -40 37288 36
rect 20456 920 37288 996
rect 20456 1880 37288 1956
rect 20456 2840 37288 2916
rect 20456 3800 37288 3876
rect 20456 4760 37288 4836
rect 20456 5720 37288 5796
rect 20456 6680 37288 6756
rect 20456 7640 37288 7716
rect 20456 8600 37288 8676
rect 20456 9560 37288 9636
rect 20456 10520 37288 10596
rect 20456 11480 37288 11556
rect 20456 12440 37288 12516
rect 20456 13400 37288 13476
rect 20456 14360 37288 14436
rect 20456 15320 37288 15396
rect 20456 16280 37288 16356
rect 20456 17240 37288 17316
rect 20456 18200 37288 18276
rect 20456 19160 37288 19236
rect 20456 20120 37288 20196
rect 20456 21080 37288 21156
rect 20456 22040 37288 22116
rect 20456 23000 37288 23076
rect 20456 23960 37288 24036
rect 20456 24920 37288 24996
rect 37288 -40 37364 24996
<< m1 >>
rect 108 7770 390 7830
rect 390 3190 2268 3250
rect 390 3190 450 7838
rect 108 16930 534 16990
rect 534 12350 2268 12410
rect 534 12350 594 16998
rect 2268 21510 2490 21570
rect 2490 3640 3796 3700
rect 2490 4600 3796 4660
rect 2490 5560 3796 5620
rect 2490 6520 3796 6580
rect 2490 7480 3796 7540
rect 2490 8440 3796 8500
rect 2490 9400 3796 9460
rect 2490 10360 3796 10420
rect 2490 11320 3796 11380
rect 2490 12280 3796 12340
rect 2490 13240 3796 13300
rect 2490 14200 3796 14260
rect 2490 15160 3796 15220
rect 2490 16120 3796 16180
rect 2490 17080 3796 17140
rect 2490 18040 3796 18100
rect 2490 19000 3796 19060
rect 2490 19960 3796 20020
rect 2490 20920 3796 20980
rect 2490 21880 3796 21940
rect 2490 22840 3796 22900
rect 2490 23800 3796 23860
rect 2490 24760 3796 24820
rect 2490 25720 3796 25780
rect 2490 3640 2550 25796
<< m2 >>
rect 108 12350 398 12426
rect 398 7770 2268 7846
rect 398 7770 474 12426
rect 108 21510 686 21586
rect 686 16930 2268 17006
rect 686 16930 762 21586
rect 108 3190 334 3266
rect 334 760 3796 836
rect 334 1720 3796 1796
rect 334 2680 3796 2756
rect 334 760 410 3266
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa10
transform 1 0 0 0 1 440
box 0 440 3656 4580
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa20
transform 1 0 0 0 1 5020
box 0 5020 3656 9160
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa30
transform 1 0 0 0 1 9600
box 0 9600 3656 13740
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa40
transform 1 0 0 0 1 14180
box 0 14180 3656 18320
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_100k xa50
transform 1 0 0 0 1 18760
box 0 18760 3656 22900
use CAP_LPF xb10
transform -1 0 37336 0 1 0
box 37336 0 71016 960
use CAP_LPF xb20
transform -1 0 37336 0 1 960
box 37336 960 71016 1920
use CAP_LPF xb21
transform -1 0 37336 0 1 1920
box 37336 1920 71016 2880
use CAP_LPF xb30
transform -1 0 37336 0 1 2880
box 37336 2880 71016 3840
use CAP_LPF xb31
transform -1 0 37336 0 1 3840
box 37336 3840 71016 4800
use CAP_LPF xb32
transform -1 0 37336 0 1 4800
box 37336 4800 71016 5760
use CAP_LPF xb33
transform -1 0 37336 0 1 5760
box 37336 5760 71016 6720
use CAP_LPF xb34
transform -1 0 37336 0 1 6720
box 37336 6720 71016 7680
use CAP_LPF xb35
transform -1 0 37336 0 1 7680
box 37336 7680 71016 8640
use CAP_LPF xb36
transform -1 0 37336 0 1 8640
box 37336 8640 71016 9600
use CAP_LPF xb37
transform -1 0 37336 0 1 9600
box 37336 9600 71016 10560
use CAP_LPF xb38
transform -1 0 37336 0 1 10560
box 37336 10560 71016 11520
use CAP_LPF xb39
transform -1 0 37336 0 1 11520
box 37336 11520 71016 12480
use CAP_LPF xb310
transform -1 0 37336 0 1 12480
box 37336 12480 71016 13440
use CAP_LPF xb311
transform -1 0 37336 0 1 13440
box 37336 13440 71016 14400
use CAP_LPF xb312
transform -1 0 37336 0 1 14400
box 37336 14400 71016 15360
use CAP_LPF xb313
transform -1 0 37336 0 1 15360
box 37336 15360 71016 16320
use CAP_LPF xb314
transform -1 0 37336 0 1 16320
box 37336 16320 71016 17280
use CAP_LPF xb315
transform -1 0 37336 0 1 17280
box 37336 17280 71016 18240
use CAP_LPF xb316
transform -1 0 37336 0 1 18240
box 37336 18240 71016 19200
use CAP_LPF xb317
transform -1 0 37336 0 1 19200
box 37336 19200 71016 20160
use CAP_LPF xb318
transform -1 0 37336 0 1 20160
box 37336 20160 71016 21120
use CAP_LPF xb319
transform -1 0 37336 0 1 21120
box 37336 21120 71016 22080
use CAP_LPF xb320
transform -1 0 37336 0 1 22080
box 37336 22080 71016 23040
use CAP_LPF xb321
transform -1 0 37336 0 1 23040
box 37336 23040 71016 24000
use CAP_LPF xb322
transform -1 0 37336 0 1 24000
box 37336 24000 71016 24960
use CAP_LPF xb323
transform -1 0 37336 0 1 24960
box 37336 24960 71016 25920
use cut_M1M4_2x1 
transform 1 0 20356 0 1 -1104
box 20356 -1104 20556 -1028
use cut_M1M2_2x1 
transform 1 0 -54 0 1 7770
box -54 7770 130 7838
use cut_M1M2_2x1 
transform 1 0 2106 0 1 3190
box 2106 3190 2290 3258
use cut_M1M3_2x1 
transform 1 0 -54 0 1 12350
box -54 12350 146 12426
use cut_M1M3_2x1 
transform 1 0 2106 0 1 7770
box 2106 7770 2306 7846
use cut_M1M2_2x1 
transform 1 0 -54 0 1 16930
box -54 16930 130 16998
use cut_M1M2_2x1 
transform 1 0 2106 0 1 12350
box 2106 12350 2290 12418
use cut_M1M3_2x1 
transform 1 0 -54 0 1 21510
box -54 21510 146 21586
use cut_M1M3_2x1 
transform 1 0 2106 0 1 16930
box 2106 16930 2306 17006
use cut_M1M2_2x1 
transform 1 0 2106 0 1 21510
box 2106 21510 2290 21578
use cut_M2M4_2x1 
transform 1 0 3696 0 1 3640
box 3696 3640 3896 3716
use cut_M2M4_2x1 
transform 1 0 3696 0 1 4600
box 3696 4600 3896 4676
use cut_M2M4_2x1 
transform 1 0 3696 0 1 5560
box 3696 5560 3896 5636
use cut_M2M4_2x1 
transform 1 0 3696 0 1 6520
box 3696 6520 3896 6596
use cut_M2M4_2x1 
transform 1 0 3696 0 1 7480
box 3696 7480 3896 7556
use cut_M2M4_2x1 
transform 1 0 3696 0 1 8440
box 3696 8440 3896 8516
use cut_M2M4_2x1 
transform 1 0 3696 0 1 9400
box 3696 9400 3896 9476
use cut_M2M4_2x1 
transform 1 0 3696 0 1 10360
box 3696 10360 3896 10436
use cut_M2M4_2x1 
transform 1 0 3696 0 1 11320
box 3696 11320 3896 11396
use cut_M2M4_2x1 
transform 1 0 3696 0 1 12280
box 3696 12280 3896 12356
use cut_M2M4_2x1 
transform 1 0 3696 0 1 13240
box 3696 13240 3896 13316
use cut_M2M4_2x1 
transform 1 0 3696 0 1 14200
box 3696 14200 3896 14276
use cut_M2M4_2x1 
transform 1 0 3696 0 1 15160
box 3696 15160 3896 15236
use cut_M2M4_2x1 
transform 1 0 3696 0 1 16120
box 3696 16120 3896 16196
use cut_M2M4_2x1 
transform 1 0 3696 0 1 17080
box 3696 17080 3896 17156
use cut_M2M4_2x1 
transform 1 0 3696 0 1 18040
box 3696 18040 3896 18116
use cut_M2M4_2x1 
transform 1 0 3696 0 1 19000
box 3696 19000 3896 19076
use cut_M2M4_2x1 
transform 1 0 3696 0 1 19960
box 3696 19960 3896 20036
use cut_M2M4_2x1 
transform 1 0 3696 0 1 20920
box 3696 20920 3896 20996
use cut_M2M4_2x1 
transform 1 0 3696 0 1 21880
box 3696 21880 3896 21956
use cut_M2M4_2x1 
transform 1 0 3696 0 1 22840
box 3696 22840 3896 22916
use cut_M2M4_2x1 
transform 1 0 3696 0 1 23800
box 3696 23800 3896 23876
use cut_M2M4_2x1 
transform 1 0 3696 0 1 24760
box 3696 24760 3896 24836
use cut_M2M4_2x1 
transform 1 0 3696 0 1 25720
box 3696 25720 3896 25796
use cut_M1M3_2x1 
transform 1 0 -54 0 1 3190
box -54 3190 146 3266
use cut_M3M4_2x1 
transform 1 0 3696 0 1 760
box 3696 760 3896 836
use cut_M3M4_2x1 
transform 1 0 3696 0 1 1720
box 3696 1720 3896 1796
use cut_M3M4_2x1 
transform 1 0 3696 0 1 2680
box 3696 2680 3896 2756
<< labels >>
flabel locali s 38200 -1104 38440 27024 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 2106 21510 2430 21730 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew
flabel locali s -54 3190 270 3410 0 FreeSans 400 0 0 0 VLPF
port 3 nsew
<< end >>
