magic
tech sky130A
magscale 1 2
timestamp 1661019234
<< checkpaint >>
rect -384 -384 1644 18336
<< locali >>
rect 1404 -384 1644 18336
rect -384 -384 1644 -144
rect -384 18096 1644 18336
rect -384 -384 -144 18336
rect 1404 -384 1644 18336
rect 432 146 600 206
rect 600 146 660 206
rect 636 294 816 354
rect 636 1994 864 2054
rect 432 498 636 558
rect 636 3754 864 3814
rect 432 2258 636 2318
rect 636 5514 864 5574
rect 432 4018 636 4078
rect 636 7274 864 7334
rect 432 5778 636 5838
rect 636 9034 864 9094
rect 432 7538 636 7598
rect 636 10794 864 10854
rect 432 9298 636 9358
rect 636 12554 864 12614
rect 432 11058 636 11118
rect 636 14314 864 14374
rect 432 12818 636 12878
rect 636 16074 864 16134
rect 432 14578 636 14638
rect 636 17834 864 17894
rect 432 16338 636 16398
rect 636 294 696 17894
rect 756 234 864 294
rect 756 234 972 294
rect 324 146 540 206
<< m3 >>
rect 756 -384 972 118
rect -108 -384 108 220
rect 756 -384 972 470
rect -108 -384 108 572
rect 756 -384 972 2230
rect -108 -384 108 2332
rect 756 -384 972 3990
rect -108 -384 108 4092
rect 756 -384 972 5750
rect -108 -384 108 5852
rect 756 -384 972 7510
rect -108 -384 108 7612
rect 756 -384 972 9270
rect -108 -384 108 9372
rect 756 -384 972 11030
rect -108 -384 108 11132
rect 756 -384 972 12790
rect -108 -384 108 12892
rect 756 -384 972 14550
rect -108 -384 108 14652
rect 756 -384 972 16310
rect -108 -384 108 16412
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa20
transform 1 0 0 0 1 0
box 0 0 1260 352
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa30
transform 1 0 0 0 1 352
box 0 352 1260 2112
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa31
transform 1 0 0 0 1 2112
box 0 2112 1260 3872
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa32
transform 1 0 0 0 1 3872
box 0 3872 1260 5632
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa33
transform 1 0 0 0 1 5632
box 0 5632 1260 7392
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa34
transform 1 0 0 0 1 7392
box 0 7392 1260 9152
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa35
transform 1 0 0 0 1 9152
box 0 9152 1260 10912
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa36
transform 1 0 0 0 1 10912
box 0 10912 1260 12672
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa37
transform 1 0 0 0 1 12672
box 0 12672 1260 14432
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa38
transform 1 0 0 0 1 14432
box 0 14432 1260 16192
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa39
transform 1 0 0 0 1 16192
box 0 16192 1260 17952
use cut_M1M4_2x1 
transform 1 0 764 0 1 58
box 764 58 964 134
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 132
box -100 132 100 208
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 410
box 764 410 964 486
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 484
box -100 484 100 560
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 2170
box 764 2170 964 2246
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 2244
box -100 2244 100 2320
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 3930
box 764 3930 964 4006
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 4004
box -100 4004 100 4080
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 5690
box 764 5690 964 5766
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 5764
box -100 5764 100 5840
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 7450
box 764 7450 964 7526
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 7524
box -100 7524 100 7600
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 9210
box 764 9210 964 9286
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 9284
box -100 9284 100 9360
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 10970
box 764 10970 964 11046
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 11044
box -100 11044 100 11120
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 12730
box 764 12730 964 12806
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 12804
box -100 12804 100 12880
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 14490
box 764 14490 964 14566
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 14564
box -100 14564 100 14640
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
use cut_M1M4_2x1 
transform 1 0 764 0 1 16250
box 764 16250 964 16326
use cut_M1M4_2x1 
transform 1 0 764 0 1 -384
box 764 -384 964 -308
use cut_M1M4_2x1 
transform 1 0 -100 0 1 16324
box -100 16324 100 16400
use cut_M1M4_2x1 
transform 1 0 -100 0 1 -384
box -100 -384 100 -308
<< labels >>
flabel locali s 1404 -384 1644 18336 0 FreeSans 400 0 0 0 AVSS
port 3 nsew
flabel locali s 756 234 972 294 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 2 nsew
<< end >>
