magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect -356 0 23524 37426
<< m3 >>
rect 8580 17456 23334 17524
rect 8580 17836 23334 17904
rect 21634 18176 21702 25396
rect 21878 18176 21946 32436
rect 4834 18284 4902 28592
rect 5550 18474 5618 28592
rect 9034 18664 9102 28592
rect 1350 18854 1418 28592
rect 1350 18854 1418 28592
rect 12738 19044 12806 28614
rect 12738 19044 12806 28614
rect 16938 19234 17006 28614
rect 16938 19234 17006 28614
rect 10362 19424 10430 28614
rect 10362 19424 10430 28614
rect 14562 19614 14630 28614
rect 14562 19614 14630 28614
rect 1962 19804 2030 28614
rect 6162 19994 6230 28614
rect 6162 19994 6230 28614
rect 4338 20184 4406 28614
rect 4338 20184 4406 28614
rect 8538 20374 8606 28614
rect 8538 20374 8606 28614
rect 2098 20564 2166 29894
rect 8402 20754 8470 29894
rect 6298 20944 6366 29894
rect 4202 21134 4270 29894
rect 10634 21324 10702 31174
rect 12466 21514 12534 31174
rect 14834 21704 14902 31174
rect 8266 21894 8334 31174
rect 4066 22084 4134 31174
rect 2234 22274 2302 31174
rect 16666 22464 16734 31174
rect 6434 22654 6502 31174
rect 10774 46 10958 114
rect 12210 46 12394 114
rect 18762 28614 18830 28798
rect 2854 27716 3038 27900
rect 8910 0 9094 4800
rect 9570 0 9754 4800
<< m2 >>
rect 14500 16954 14568 17524
rect 8580 16954 8648 17904
rect 4834 18216 13624 18284
rect 5550 18406 13248 18474
rect 9034 18596 12872 18664
rect 1350 18786 14000 18854
rect 10848 18976 12806 19044
rect 11224 19166 17006 19234
rect 10362 19356 10728 19424
rect 11036 19546 14630 19614
rect 1962 19736 9224 19804
rect 6162 19926 9976 19994
rect 4338 20116 9600 20184
rect 8538 20306 10352 20374
rect 2098 20496 9412 20564
rect 8402 20686 10540 20754
rect 6298 20876 10164 20944
rect 4202 21066 9788 21134
rect 10634 21256 12496 21324
rect 12240 21446 12534 21514
rect 12052 21636 14902 21704
rect 8266 21826 12684 21894
rect 4066 22016 13436 22084
rect 2234 22206 13812 22274
rect 11864 22396 16734 22464
rect 6434 22586 13060 22654
rect 1350 23792 1534 23860
<< m4 >>
rect 21634 17836 21702 18176
rect 21878 17456 21946 18176
<< m1 >>
rect 13556 16894 13624 18216
rect 13180 16894 13248 18406
rect 12804 16894 12872 18596
rect 13932 16894 14000 18786
rect 10848 16894 10916 18976
rect 11224 16894 11292 19166
rect 10660 16894 10728 19356
rect 11036 16894 11104 19546
rect 9156 16894 9224 19736
rect 9908 16894 9976 19926
rect 9532 16894 9600 20116
rect 10284 16894 10352 20306
rect 9344 16894 9412 20496
rect 10472 16894 10540 20686
rect 10096 16894 10164 20876
rect 9720 16894 9788 21066
rect 12428 16894 12496 21256
rect 12240 16894 12308 21446
rect 12052 16894 12120 21636
rect 12616 16894 12684 21826
rect 13368 16894 13436 22016
rect 13744 16894 13812 22206
rect 11864 16894 11932 22396
rect 12992 16894 13060 22586
<< locali >>
rect 10774 2450 10954 2510
rect 10774 1170 10954 1230
rect 18514 34116 18694 34176
rect 1354 32756 1534 32816
rect 9934 450 10114 510
use SARBSSW_CV XB1
transform -1 0 11584 0 1 0
box 11584 0 23524 4800
use SARBSSW_CV XB2
transform 1 0 11584 0 1 0
box 11584 0 23524 4800
use CDAC8_CV XDAC1
transform -1 0 11404 0 1 4990
box 11404 4990 22692 16954
use CDAC8_CV XDAC2
transform 1 0 11744 0 1 4990
box 11744 4990 23032 16954
use SARDIGEX4_CV XA0
transform 1 0 1084 0 1 23346
box 1084 23346 3184 36466
use SARDIGEX4_CV XA1
transform -1 0 5284 0 1 23346
box 5284 23346 7384 36466
use SARDIGEX4_CV XA2
transform 1 0 5284 0 1 23346
box 5284 23346 7384 36466
use SARDIGEX4_CV XA3
transform -1 0 9484 0 1 23346
box 9484 23346 11584 36466
use SARDIGEX4_CV XA4
transform 1 0 9484 0 1 23346
box 9484 23346 11584 36466
use SARDIGEX4_CV XA5
transform -1 0 13684 0 1 23346
box 13684 23346 15784 36466
use SARDIGEX4_CV XA6
transform 1 0 13684 0 1 23346
box 13684 23346 15784 36466
use SARDIGEX4_CV XA7
transform -1 0 17884 0 1 23346
box 17884 23346 19984 36466
use SARDIGEX4_CV XA8
transform 1 0 17884 0 1 23346
box 17884 23346 19984 36466
use SARCMPX1_CV XA20
transform -1 0 22084 0 1 23346
box 22084 23346 24184 37426
use cut_M3M4_1x2 
transform 1 0 14500 0 1 16954
box 14500 16954 14568 17138
use cut_M3M4_2x1 
transform 1 0 14500 0 1 17456
box 14500 17456 14684 17524
use cut_M3M4_1x2 
transform 1 0 8580 0 1 16954
box 8580 16954 8648 17138
use cut_M3M4_2x1 
transform 1 0 8580 0 1 17836
box 8580 17836 8764 17904
use cut_M2M4_2x1 
transform 1 0 21634 0 1 25396
box 21634 25396 21818 25464
use cut_M4M5_2x1 
transform 1 0 21634 0 1 17836
box 21634 17836 21818 17904
use cut_M4M5_1x2 
transform 1 0 21634 0 1 18176
box 21634 18176 21702 18360
use cut_M3M4_2x1 
transform 1 0 21762 0 1 32436
box 21762 32436 21946 32504
use cut_M2M3_2x1 
transform 1 0 21634 0 1 32436
box 21634 32436 21818 32504
use cut_M4M5_2x1 
transform 1 0 21878 0 1 17456
box 21878 17456 22062 17524
use cut_M4M5_1x2 
transform 1 0 21878 0 1 18176
box 21878 18176 21946 18360
use cut_M3M4_1x2 
transform 1 0 4834 0 1 18158
box 4834 18158 4902 18342
use cut_M2M3_1x2 
transform 1 0 13552 0 1 18158
box 13552 18158 13620 18342
use cut_M3M4_1x2 
transform 1 0 5550 0 1 18348
box 5550 18348 5618 18532
use cut_M2M3_1x2 
transform 1 0 13176 0 1 18348
box 13176 18348 13244 18532
use cut_M3M4_1x2 
transform 1 0 9034 0 1 18538
box 9034 18538 9102 18722
use cut_M2M3_1x2 
transform 1 0 12800 0 1 18538
box 12800 18538 12868 18722
use cut_M3M4_1x2 
transform 1 0 1350 0 1 18728
box 1350 18728 1418 18912
use cut_M2M3_1x2 
transform 1 0 13928 0 1 18728
box 13928 18728 13996 18912
use cut_M3M4_1x2 
transform 1 0 12738 0 1 18918
box 12738 18918 12806 19102
use cut_M2M3_1x2 
transform 1 0 10844 0 1 18918
box 10844 18918 10912 19102
use cut_M3M4_1x2 
transform 1 0 16938 0 1 19108
box 16938 19108 17006 19292
use cut_M2M3_1x2 
transform 1 0 11220 0 1 19108
box 11220 19108 11288 19292
use cut_M3M4_1x2 
transform 1 0 10362 0 1 19298
box 10362 19298 10430 19482
use cut_M2M3_1x2 
transform 1 0 10656 0 1 19298
box 10656 19298 10724 19482
use cut_M3M4_1x2 
transform 1 0 14562 0 1 19488
box 14562 19488 14630 19672
use cut_M2M3_1x2 
transform 1 0 11032 0 1 19488
box 11032 19488 11100 19672
use cut_M3M4_1x2 
transform 1 0 1962 0 1 19678
box 1962 19678 2030 19862
use cut_M2M3_1x2 
transform 1 0 9152 0 1 19678
box 9152 19678 9220 19862
use cut_M3M4_1x2 
transform 1 0 6162 0 1 19868
box 6162 19868 6230 20052
use cut_M2M3_1x2 
transform 1 0 9904 0 1 19868
box 9904 19868 9972 20052
use cut_M3M4_1x2 
transform 1 0 4338 0 1 20058
box 4338 20058 4406 20242
use cut_M2M3_1x2 
transform 1 0 9528 0 1 20058
box 9528 20058 9596 20242
use cut_M3M4_1x2 
transform 1 0 8538 0 1 20248
box 8538 20248 8606 20432
use cut_M2M3_1x2 
transform 1 0 10280 0 1 20248
box 10280 20248 10348 20432
use cut_M3M4_1x2 
transform 1 0 2098 0 1 20438
box 2098 20438 2166 20622
use cut_M2M3_1x2 
transform 1 0 9340 0 1 20438
box 9340 20438 9408 20622
use cut_M3M4_1x2 
transform 1 0 8402 0 1 20628
box 8402 20628 8470 20812
use cut_M2M3_1x2 
transform 1 0 10468 0 1 20628
box 10468 20628 10536 20812
use cut_M3M4_1x2 
transform 1 0 6298 0 1 20818
box 6298 20818 6366 21002
use cut_M2M3_1x2 
transform 1 0 10092 0 1 20818
box 10092 20818 10160 21002
use cut_M3M4_1x2 
transform 1 0 4202 0 1 21008
box 4202 21008 4270 21192
use cut_M2M3_1x2 
transform 1 0 9716 0 1 21008
box 9716 21008 9784 21192
use cut_M3M4_1x2 
transform 1 0 10634 0 1 21198
box 10634 21198 10702 21382
use cut_M2M3_1x2 
transform 1 0 12424 0 1 21198
box 12424 21198 12492 21382
use cut_M3M4_1x2 
transform 1 0 12466 0 1 21388
box 12466 21388 12534 21572
use cut_M2M3_1x2 
transform 1 0 12236 0 1 21388
box 12236 21388 12304 21572
use cut_M3M4_1x2 
transform 1 0 14834 0 1 21578
box 14834 21578 14902 21762
use cut_M2M3_1x2 
transform 1 0 12048 0 1 21578
box 12048 21578 12116 21762
use cut_M3M4_1x2 
transform 1 0 8266 0 1 21768
box 8266 21768 8334 21952
use cut_M2M3_1x2 
transform 1 0 12612 0 1 21768
box 12612 21768 12680 21952
use cut_M3M4_1x2 
transform 1 0 4066 0 1 21958
box 4066 21958 4134 22142
use cut_M2M3_1x2 
transform 1 0 13364 0 1 21958
box 13364 21958 13432 22142
use cut_M3M4_1x2 
transform 1 0 2234 0 1 22148
box 2234 22148 2302 22332
use cut_M2M3_1x2 
transform 1 0 13740 0 1 22148
box 13740 22148 13808 22332
use cut_M3M4_1x2 
transform 1 0 16666 0 1 22338
box 16666 22338 16734 22522
use cut_M2M3_1x2 
transform 1 0 11860 0 1 22338
box 11860 22338 11928 22522
use cut_M3M4_1x2 
transform 1 0 6434 0 1 22528
box 6434 22528 6502 22712
use cut_M2M3_1x2 
transform 1 0 12988 0 1 22528
box 12988 22528 13056 22712
<< labels >>
flabel m3 s 1350 18854 1418 28592 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 12738 19044 12806 28614 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 16938 19234 17006 28614 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 10362 19424 10430 28614 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 14562 19614 14630 28614 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 6162 19994 6230 28614 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 4338 20184 4406 28614 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8538 20374 8606 28614 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel m3 s 10774 46 10958 114 0 FreeSans 400 0 0 0 SAR_IP
port 9 nsew
flabel m3 s 12210 46 12394 114 0 FreeSans 400 0 0 0 SAR_IN
port 10 nsew
flabel locali s 10774 2450 10954 2510 0 FreeSans 400 0 0 0 SARN
port 11 nsew
flabel locali s 10774 1170 10954 1230 0 FreeSans 400 0 0 0 SARP
port 12 nsew
flabel locali s 18514 34116 18694 34176 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 18762 28614 18830 28798 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
flabel m2 s 1350 23792 1534 23860 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s 1354 32756 1534 32816 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 9934 450 10114 510 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel m3 s 2854 27716 3038 27900 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel m3 s 8910 0 9094 4800 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel m3 s 9570 0 9754 4800 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
<< end >>
