magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 2240
<< locali >>
rect 770 210 830 2030
rect 800 210 968 270
rect 968 50 1520 110
rect 968 50 1028 270
rect 370 450 430 1790
rect 1890 450 1950 2110
rect 1490 210 1550 2190
rect 680 2130 1640 2190
rect 1520 2130 1688 2190
rect 1688 2050 1920 2110
rect 1688 2050 1748 2190
rect 770 210 830 430
rect 770 530 830 750
rect 770 850 830 1070
rect 770 1170 830 1390
rect 770 1490 830 1710
rect 770 1810 830 2030
rect 1490 210 1550 430
rect 1490 530 1550 750
rect 1490 850 1550 1070
rect 1490 1170 1550 1390
rect 1490 1490 1550 1710
rect 1490 1810 1550 2030
<< poly >>
rect 280 142 2040 178
<< m3 >>
rect 1400 0 1600 2240
rect 680 0 880 2240
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1160 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1160 1280
use NCHDL MN4
transform 1 0 0 0 1 1280
box 0 1280 1160 1600
use NCHDL MN5
transform 1 0 0 0 1 1600
box 0 1600 1160 1920
use NCHDL MN6
transform 1 0 0 0 1 1920
box 0 1920 1160 2240
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1_DMY
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL MP2_DMY
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use PCHDL MP3_DMY
transform 1 0 1160 0 1 960
box 1160 960 2320 1280
use PCHDL MP4_DMY
transform 1 0 1160 0 1 1280
box 1160 1280 2320 1600
use PCHDL MP5_DMY
transform 1 0 1160 0 1 1600
box 1160 1600 2320 1920
use PCHDL MP6_DMY
transform 1 0 1160 0 1 1920
box 1160 1920 2320 2240
use cut_M1M4_2x1 
transform 1 0 1400 0 1 210
box 1400 210 1600 278
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
<< labels >>
flabel locali s 2200 120 2440 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -120 120 120 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 280 2050 520 2110 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 CKN
port 4 nsew
flabel locali s 280 450 520 510 0 FreeSans 400 0 0 0 CI
port 5 nsew
flabel m3 s 1400 0 1600 2240 0 FreeSans 400 0 0 0 AVDD
port 6 nsew
flabel m3 s 680 0 880 2240 0 FreeSans 400 0 0 0 AVSS
port 7 nsew
<< end >>
