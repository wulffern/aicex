magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 184 68
<< m1 >>
rect 0 0 184 68
<< m2 >>
rect 0 0 184 68
<< m3 >>
rect 0 0 184 68
<< v1 >>
rect 12 6 172 62
<< v2 >>
rect 12 6 172 62
<< labels >>
<< end >>
