magic
tech sky130A
magscale 1 2
timestamp 1658775803
<< checkpaint >>
rect 0 30 984 606
<< m4 >>
rect 0 0 984 76
rect 264 140 492 216
rect 644 140 720 216
rect 0 280 984 356
rect 264 420 492 496
rect 644 420 720 496
rect 0 560 984 636
rect 0 0 76 560
rect 908 0 984 560
use cut_M4M5_2x1 
transform 1 0 64 0 1 140
box 64 140 264 216
use cut_M4M5_2x1 
transform 1 0 720 0 1 140
box 720 140 920 216
use cut_M4M5_2x1 
transform 1 0 64 0 1 420
box 64 420 264 496
use cut_M4M5_2x1 
transform 1 0 720 0 1 420
box 720 420 920 496
<< labels >>
<< end >>
