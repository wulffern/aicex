magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 1980 14080
<< locali >>
rect 1260 4530 1398 4590
rect 1398 8770 1620 8830
rect 1398 6210 1620 6270
rect 1398 4530 1458 8830
rect 162 2370 360 2430
rect 162 2690 360 2750
rect 162 7490 360 7550
rect 162 11650 360 11710
rect 162 2370 222 11710
rect 360 11650 498 11710
rect 498 12050 720 12110
rect 498 11650 558 12110
rect 522 13170 720 13230
rect 360 12290 522 12350
rect 522 12290 582 13230
rect 1260 13650 1398 13710
rect 1398 12610 1620 12670
rect 1398 12610 1458 13710
rect 522 4050 720 4110
rect 522 8850 720 8910
rect 522 4050 582 8910
<< m1 >>
rect 1260 8690 1398 8750
rect 1398 4290 1620 4350
rect 1398 4930 1620 4990
rect 1398 4290 1458 8758
rect 360 2050 498 2110
rect 360 3010 498 3070
rect 498 2050 558 3078
rect 360 9090 498 9150
rect 360 10050 498 10110
rect 498 9090 558 10118
rect 162 450 360 510
rect 162 9730 360 9790
rect 162 11970 360 12030
rect 162 450 222 12038
rect 360 11970 498 12030
rect 498 12690 720 12750
rect 498 11970 558 12758
<< m3 >>
rect 1170 0 1354 14080
rect 630 0 814 14080
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use TAPCELLB_CV XA0
transform 1 0 0 0 1 0
box 0 0 1980 320
use SARKICKHX1_CV XA1
transform 1 0 0 0 1 320
box 0 320 1980 2560
use SARCMPHX1_CV XA2
transform 1 0 0 0 1 2560
box 0 2560 1980 4800
use IVX4_CV XA2a
transform 1 0 0 0 1 4800
box 0 4800 1980 6080
use IVX4_CV XA3a
transform 1 0 0 0 1 6080
box 0 6080 1980 7360
use SARCMPHX1_CV XA3
transform 1 0 0 0 1 7360
box 0 7360 1980 9600
use SARKICKHX1_CV XA4
transform 1 0 0 0 1 9600
box 0 9600 1980 11840
use IVX1_CV XA9
transform 1 0 0 0 1 11840
box 0 11840 1980 12160
use NDX1_CV XA10
transform 1 0 0 0 1 12160
box 0 12160 1980 12800
use NRX1_CV XA11
transform 1 0 0 0 1 12800
box 0 12800 1980 13440
use IVX1_CV XA12
transform 1 0 0 0 1 13440
box 0 13440 1980 13760
use TAPCELLB_CV XA13
transform 1 0 0 0 1 13760
box 0 13760 1980 14080
use DMY_CV XA14
transform 1 0 0 0 1 14080
box 0 14080 0 14080
use cut_M1M2_2x1 
transform 1 0 1170 0 1 8690
box 1170 8690 1354 8758
use cut_M1M2_2x1 
transform 1 0 1530 0 1 4290
box 1530 4290 1714 4358
use cut_M1M2_2x1 
transform 1 0 1530 0 1 4930
box 1530 4930 1714 4998
use cut_M1M2_2x1 
transform 1 0 266 0 1 2050
box 266 2050 450 2118
use cut_M1M2_2x1 
transform 1 0 266 0 1 3010
box 266 3010 450 3078
use cut_M1M2_2x1 
transform 1 0 266 0 1 9090
box 266 9090 450 9158
use cut_M1M2_2x1 
transform 1 0 266 0 1 10050
box 266 10050 450 10118
use cut_M1M2_2x1 
transform 1 0 270 0 1 450
box 270 450 454 518
use cut_M1M2_2x1 
transform 1 0 270 0 1 9730
box 270 9730 454 9798
use cut_M1M2_2x1 
transform 1 0 270 0 1 11970
box 270 11970 454 12038
use cut_M1M2_2x1 
transform 1 0 270 0 1 11970
box 270 11970 454 12038
use cut_M1M2_2x1 
transform 1 0 630 0 1 12690
box 630 12690 814 12758
<< labels >>
flabel locali s 270 12930 450 12990 0 FreeSans 400 0 0 0 CK_SAMPLE
port 1 nsew
flabel locali s 270 13570 450 13630 0 FreeSans 400 0 0 0 CK_CMP
port 2 nsew
flabel locali s 270 13250 450 13310 0 FreeSans 400 0 0 0 DONE
port 3 nsew
flabel locali s 630 6290 810 6350 0 FreeSans 400 0 0 0 CNO
port 4 nsew
flabel locali s 630 5010 810 5070 0 FreeSans 400 0 0 0 CPO
port 5 nsew
flabel locali s 270 2050 450 2110 0 FreeSans 400 0 0 0 CPI
port 6 nsew
flabel locali s 270 9090 450 9150 0 FreeSans 400 0 0 0 CNI
port 7 nsew
flabel m3 s 1170 0 1354 14080 0 FreeSans 400 0 0 0 AVDD
port 8 nsew
flabel m3 s 630 0 814 14080 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
<< end >>
