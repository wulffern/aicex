magic
tech sky130A
magscale 1 2
timestamp 1658775803
<< checkpaint >>
rect 0 30 9504 3510
<< m3 >>
rect 328 0 404 3540
rect 328 0 404 3540
rect 468 140 544 3400
rect 608 0 684 3540
rect 748 140 824 3400
rect 888 0 964 3540
rect 1028 140 1104 3400
rect 1168 0 1244 3540
rect 1308 140 1384 3400
rect 1448 0 1524 3540
rect 1588 140 1664 3400
rect 1728 0 1804 3540
rect 1868 140 1944 3400
rect 2008 0 2084 3540
rect 2148 140 2224 3400
rect 2288 0 2364 3540
rect 2428 140 2504 3400
rect 2568 0 2644 3540
rect 2708 140 2784 3400
rect 2848 0 2924 3540
rect 2988 140 3064 3400
rect 3128 0 3204 3540
rect 3268 140 3344 3400
rect 3408 0 3484 3540
rect 3548 140 3624 3400
rect 3688 0 3764 3540
rect 3828 140 3904 3400
rect 3968 0 4044 3540
rect 4108 140 4184 3400
rect 4248 0 4324 3540
rect 4388 140 4464 3400
rect 4528 0 4604 3540
rect 4668 140 4744 3400
rect 4808 0 4884 3540
rect 4948 140 5024 3400
rect 5088 0 5164 3540
rect 5228 140 5304 3400
rect 5368 0 5444 3540
rect 5508 140 5584 3400
rect 5648 0 5724 3540
rect 5788 140 5864 3400
rect 5928 0 6004 3540
rect 6068 140 6144 3400
rect 6208 0 6284 3540
rect 6348 140 6424 3400
rect 6488 0 6564 3540
rect 6628 140 6704 3400
rect 6768 0 6844 3540
rect 6908 140 6984 3400
rect 7048 0 7124 3540
rect 7188 140 7264 3400
rect 7328 0 7404 3540
rect 7468 140 7544 3400
rect 7608 0 7684 3540
rect 7748 140 7824 3400
rect 7888 0 7964 3540
rect 8028 140 8104 3400
rect 8168 0 8244 3540
rect 8308 140 8384 3400
rect 8448 0 8524 3540
rect 8588 140 8664 3400
rect 8728 0 8804 3540
rect 8868 140 8944 3400
rect 9008 0 9084 3540
rect 9148 140 9224 3400
rect 9428 0 9504 3540
rect 9288 0 9364 3540
rect 328 0 9288 76
rect 328 3464 9288 3540
<< m1 >>
rect 328 0 9428 76
rect 2428 400 2504 3540
rect 7188 0 7264 3140
rect 2708 0 2784 1304
rect 2708 1624 2784 3540
rect 6908 0 6984 1304
rect 6908 1624 6984 3540
rect 2148 0 2224 2528
rect 2148 2848 2224 3540
rect 2988 0 3064 2528
rect 2988 2848 3064 3540
rect 6628 0 6704 2528
rect 6628 2848 6704 3540
rect 7468 0 7544 2528
rect 7468 2848 7544 3540
rect 1588 0 1664 1916
rect 1588 2236 1664 3540
rect 1868 0 1944 1916
rect 1868 2236 1944 3540
rect 3268 0 3344 1916
rect 3268 2236 3344 3540
rect 3548 0 3624 1916
rect 3548 2236 3624 3540
rect 6068 0 6144 1916
rect 6068 2236 6144 3540
rect 6348 0 6424 1916
rect 6348 2236 6424 3540
rect 7748 0 7824 1916
rect 7748 2236 7824 3540
rect 8028 0 8104 1916
rect 8028 2236 8104 3540
rect 468 0 544 692
rect 468 1012 544 3540
rect 748 0 824 692
rect 748 1012 824 3540
rect 1028 0 1104 692
rect 1028 1012 1104 3540
rect 1308 0 1384 692
rect 1308 1012 1384 3540
rect 3828 0 3904 692
rect 3828 1012 3904 3540
rect 4108 0 4184 692
rect 4108 1012 4184 3540
rect 4388 0 4464 692
rect 4388 1012 4464 3540
rect 4668 0 4744 692
rect 4668 1012 4744 3540
rect 4948 0 5024 692
rect 4948 1012 5024 3540
rect 5228 0 5304 692
rect 5228 1012 5304 3540
rect 5508 0 5584 692
rect 5508 1012 5584 3540
rect 5788 0 5864 692
rect 5788 1012 5864 3540
rect 8308 0 8384 692
rect 8308 1012 8384 3540
rect 8588 0 8664 692
rect 8588 1012 8664 3540
rect 8868 0 8944 692
rect 8868 1012 8944 3540
rect 9148 0 9224 692
rect 9148 1012 9224 3540
rect 328 0 404 3464
rect 608 0 684 3464
rect 888 0 964 3464
rect 1168 0 1244 3464
rect 1448 0 1524 3464
rect 1728 0 1804 3464
rect 2008 0 2084 3464
rect 2288 0 2364 3464
rect 2568 0 2644 3464
rect 2848 0 2924 3464
rect 3128 0 3204 3464
rect 3408 0 3484 3464
rect 3688 0 3764 3464
rect 3968 0 4044 3464
rect 4248 0 4324 3464
rect 4528 0 4604 3464
rect 4808 0 4884 3464
rect 5088 0 5164 3464
rect 5368 0 5444 3464
rect 5648 0 5724 3464
rect 5928 0 6004 3464
rect 6208 0 6284 3464
rect 6488 0 6564 3464
rect 6768 0 6844 3464
rect 7048 0 7124 3464
rect 7328 0 7404 3464
rect 7608 0 7684 3464
rect 7888 0 7964 3464
rect 8168 0 8244 3464
rect 8448 0 8524 3464
rect 8728 0 8804 3464
rect 9008 0 9084 3464
rect 9428 0 9504 3540
rect 9288 0 9364 3540
rect 328 0 9428 76
rect 328 3464 9428 3540
<< locali >>
rect 0 202 200 278
rect 0 3262 200 3338
rect 0 1426 200 1502
rect 0 2650 200 2726
rect 0 2038 200 2114
rect 0 814 200 890
rect 320 814 9288 890
rect 320 202 9288 278
rect 320 3262 9288 3338
rect 320 1426 9288 1502
rect 320 2650 9288 2726
rect 320 2038 9288 2114
<< m4 >>
rect 188 0 264 3540
rect 468 0 544 3540
rect 748 0 824 3540
rect 1028 0 1104 3540
rect 1308 0 1384 3540
rect 1588 0 1664 3540
rect 1868 0 1944 3540
rect 2148 0 2224 3540
rect 2428 0 2504 3540
rect 2708 0 2784 3540
rect 2988 0 3064 3540
rect 3268 0 3344 3540
rect 3548 0 3624 3540
rect 3828 0 3904 3540
rect 4108 0 4184 3540
rect 4388 0 4464 3540
rect 4668 0 4744 3540
rect 4948 0 5024 3540
rect 5228 0 5304 3540
rect 5508 0 5584 3540
rect 5788 0 5864 3540
rect 6068 0 6144 3540
rect 6348 0 6424 3540
rect 6628 0 6704 3540
rect 6908 0 6984 3540
rect 7188 0 7264 3540
rect 7468 0 7544 3540
rect 7748 0 7824 3540
rect 8028 0 8104 3540
rect 8308 0 8384 3540
rect 8588 0 8664 3540
rect 8868 0 8944 3540
rect 9148 0 9224 3540
rect 9428 0 9504 3540
rect 188 0 9428 76
rect 188 3464 9428 3540
<< m2 >>
rect 9428 0 9504 3540
use RM1 XRES1A
transform 1 0 200 0 1 202
box 200 202 320 202
use RM1 XRES1B
transform 1 0 200 0 1 3262
box 200 3262 320 3262
use RM1 XRES2
transform 1 0 200 0 1 1426
box 200 1426 320 1426
use RM1 XRES4
transform 1 0 200 0 1 2650
box 200 2650 320 2650
use RM1 XRES8
transform 1 0 200 0 1 2038
box 200 2038 320 2038
use RM1 XRES16
transform 1 0 200 0 1 814
box 200 814 320 814
use cut_M2M5_1x2 
transform 1 0 9428 0 1 1570
box 9428 1570 9504 1770
use cut_M1M4_1x2 
transform 1 0 2428 0 1 140
box 2428 140 2504 340
use cut_M1M4_1x2 
transform 1 0 7188 0 1 3200
box 7188 3200 7264 3400
use cut_M1M4_1x2 
transform 1 0 2708 0 1 1364
box 2708 1364 2784 1564
use cut_M1M4_1x2 
transform 1 0 6908 0 1 1364
box 6908 1364 6984 1564
use cut_M1M4_1x2 
transform 1 0 2148 0 1 2588
box 2148 2588 2224 2788
use cut_M1M4_1x2 
transform 1 0 2988 0 1 2588
box 2988 2588 3064 2788
use cut_M1M4_1x2 
transform 1 0 6628 0 1 2588
box 6628 2588 6704 2788
use cut_M1M4_1x2 
transform 1 0 7468 0 1 2588
box 7468 2588 7544 2788
use cut_M1M4_1x2 
transform 1 0 1588 0 1 1976
box 1588 1976 1664 2176
use cut_M1M4_1x2 
transform 1 0 1868 0 1 1976
box 1868 1976 1944 2176
use cut_M1M4_1x2 
transform 1 0 3268 0 1 1976
box 3268 1976 3344 2176
use cut_M1M4_1x2 
transform 1 0 3548 0 1 1976
box 3548 1976 3624 2176
use cut_M1M4_1x2 
transform 1 0 6068 0 1 1976
box 6068 1976 6144 2176
use cut_M1M4_1x2 
transform 1 0 6348 0 1 1976
box 6348 1976 6424 2176
use cut_M1M4_1x2 
transform 1 0 7748 0 1 1976
box 7748 1976 7824 2176
use cut_M1M4_1x2 
transform 1 0 8028 0 1 1976
box 8028 1976 8104 2176
use cut_M1M4_1x2 
transform 1 0 468 0 1 752
box 468 752 544 952
use cut_M1M4_1x2 
transform 1 0 748 0 1 752
box 748 752 824 952
use cut_M1M4_1x2 
transform 1 0 1028 0 1 752
box 1028 752 1104 952
use cut_M1M4_1x2 
transform 1 0 1308 0 1 752
box 1308 752 1384 952
use cut_M1M4_1x2 
transform 1 0 3828 0 1 752
box 3828 752 3904 952
use cut_M1M4_1x2 
transform 1 0 4108 0 1 752
box 4108 752 4184 952
use cut_M1M4_1x2 
transform 1 0 4388 0 1 752
box 4388 752 4464 952
use cut_M1M4_1x2 
transform 1 0 4668 0 1 752
box 4668 752 4744 952
use cut_M1M4_1x2 
transform 1 0 4948 0 1 752
box 4948 752 5024 952
use cut_M1M4_1x2 
transform 1 0 5228 0 1 752
box 5228 752 5304 952
use cut_M1M4_1x2 
transform 1 0 5508 0 1 752
box 5508 752 5584 952
use cut_M1M4_1x2 
transform 1 0 5788 0 1 752
box 5788 752 5864 952
use cut_M1M4_1x2 
transform 1 0 8308 0 1 752
box 8308 752 8384 952
use cut_M1M4_1x2 
transform 1 0 8588 0 1 752
box 8588 752 8664 952
use cut_M1M4_1x2 
transform 1 0 8868 0 1 752
box 8868 752 8944 952
use cut_M1M4_1x2 
transform 1 0 9148 0 1 752
box 9148 752 9224 952
<< labels >>
flabel m3 s 328 0 404 3540 0 FreeSans 400 0 0 0 CTOP
port 7 nsew
flabel m1 s 328 0 9428 76 0 FreeSans 400 0 0 0 AVSS
port 8 nsew
flabel locali s 0 202 200 278 0 FreeSans 400 0 0 0 C1A
port 1 nsew
flabel locali s 0 3262 200 3338 0 FreeSans 400 0 0 0 C1B
port 2 nsew
flabel locali s 0 1426 200 1502 0 FreeSans 400 0 0 0 C2
port 3 nsew
flabel locali s 0 2650 200 2726 0 FreeSans 400 0 0 0 C4
port 4 nsew
flabel locali s 0 2038 200 2114 0 FreeSans 400 0 0 0 C8
port 5 nsew
flabel locali s 0 814 200 890 0 FreeSans 400 0 0 0 C16
port 6 nsew
<< end >>
