magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect -4072 0 26328 37462
<< m3 >>
rect 8580 17864 26150 17924
rect 8580 18220 26150 18280
rect 22208 18552 22268 25432
rect 22496 18552 22556 32472
rect 3648 18636 3708 28628
rect 4488 18814 4548 28628
rect 8288 18992 8348 28628
rect -152 19170 -92 28628
rect 12324 19348 12384 28642
rect 16964 19526 17024 28642
rect 9864 19704 9924 28642
rect 14504 19882 14564 28642
rect 584 20060 644 28642
rect 5224 20238 5284 28642
rect 3044 20416 3104 28642
rect 7684 20594 7744 28642
rect 720 20772 780 29922
rect 7548 20950 7608 29922
rect 5360 21128 5420 29922
rect 2908 21306 2968 29922
rect 10136 21484 10196 31202
rect 12052 21662 12112 31202
rect 14776 21840 14836 31202
rect 7412 22018 7472 31202
rect 2772 22196 2832 31202
rect 856 22374 916 31202
rect 16692 22552 16752 31202
rect 5496 22730 5556 31202
<< m2 >>
rect 13604 17390 13664 17932
rect 8580 17390 8640 18288
rect 3648 18576 12832 18636
rect 4488 18754 12520 18814
rect 8288 18932 12208 18992
rect -152 19110 13144 19170
rect 10512 19288 12384 19348
rect 10824 19466 17024 19526
rect 9864 19644 10416 19704
rect 10668 19822 14564 19882
rect 584 20000 9168 20060
rect 5224 20178 9792 20238
rect 3044 20356 9480 20416
rect 7684 20534 10104 20594
rect 720 20712 9324 20772
rect 7548 20890 10260 20950
rect 5360 21068 9948 21128
rect 2908 21246 9636 21306
rect 10136 21424 11896 21484
rect 11680 21602 12112 21662
rect 11524 21780 14836 21840
rect 7412 21958 12052 22018
rect 2772 22136 12676 22196
rect 856 22314 12988 22374
rect 11368 22492 16752 22552
rect 5496 22670 12364 22730
<< m4 >>
rect 22208 18220 22268 18552
rect 22496 17864 22556 18552
<< m1 >>
rect 12772 17330 12832 18576
rect 12460 17330 12520 18754
rect 12148 17330 12208 18932
rect 13084 17330 13144 19110
rect 10512 17330 10572 19288
rect 10824 17330 10884 19466
rect 10356 17330 10416 19644
rect 10668 17330 10728 19822
rect 9108 17330 9168 20000
rect 9732 17330 9792 20178
rect 9420 17330 9480 20356
rect 10044 17330 10104 20534
rect 9264 17330 9324 20712
rect 10200 17330 10260 20890
rect 9888 17330 9948 21068
rect 9576 17330 9636 21246
rect 11836 17330 11896 21424
rect 11680 17330 11740 21602
rect 11524 17330 11584 21780
rect 11992 17330 12052 21958
rect 12616 17330 12676 22136
rect 12928 17330 12988 22314
rect 11368 17330 11428 22492
rect 12304 17330 12364 22670
use SARBSSW_CV XB1
transform -1 0 11128 0 1 0
box 11128 0 26328 4800
use SARBSSW_CV XB2
transform 1 0 11128 0 1 0
box 11128 0 26328 4800
use CDAC8_CV XDAC1
transform -1 0 11004 0 1 4978
box 11004 4978 21892 17390
use CDAC8_CV XDAC2
transform 1 0 11248 0 1 4978
box 11248 4978 22136 17390
use SARDIGEX4_CV XA0
transform 1 0 -472 0 1 23382
box -472 23382 1848 36502
use SARDIGEX4_CV XA1
transform -1 0 4168 0 1 23382
box 4168 23382 6488 36502
use SARDIGEX4_CV XA2
transform 1 0 4168 0 1 23382
box 4168 23382 6488 36502
use SARDIGEX4_CV XA3
transform -1 0 8808 0 1 23382
box 8808 23382 11128 36502
use SARDIGEX4_CV XA4
transform 1 0 8808 0 1 23382
box 8808 23382 11128 36502
use SARDIGEX4_CV XA5
transform -1 0 13448 0 1 23382
box 13448 23382 15768 36502
use SARDIGEX4_CV XA6
transform 1 0 13448 0 1 23382
box 13448 23382 15768 36502
use SARDIGEX4_CV XA7
transform -1 0 18088 0 1 23382
box 18088 23382 20408 36502
use SARDIGEX4_CV XA8
transform 1 0 18088 0 1 23382
box 18088 23382 20408 36502
use SARCMPX1_CV XA20
transform -1 0 22728 0 1 23382
box 22728 23382 25048 37462
use cut_M3M4_1x2 
transform 1 0 13604 0 1 17390
box 13604 17390 13672 17590
use cut_M3M4_2x1 
transform 1 0 13604 0 1 17864
box 13604 17864 13804 17932
use cut_M3M4_1x2 
transform 1 0 8580 0 1 17390
box 8580 17390 8648 17590
use cut_M3M4_2x1 
transform 1 0 8580 0 1 18220
box 8580 18220 8780 18288
use cut_M2M4_2x1 
transform 1 0 22208 0 1 25432
box 22208 25432 22408 25500
use cut_M4M5_2x1 
transform 1 0 22208 0 1 18220
box 22208 18220 22408 18288
use cut_M4M5_1x2 
transform 1 0 22208 0 1 18552
box 22208 18552 22276 18752
use cut_M3M4_2x1 
transform 1 0 22356 0 1 32472
box 22356 32472 22556 32540
use cut_M2M3_2x1 
transform 1 0 22208 0 1 32472
box 22208 32472 22408 32540
use cut_M4M5_2x1 
transform 1 0 22496 0 1 17864
box 22496 17864 22696 17932
use cut_M4M5_1x2 
transform 1 0 22496 0 1 18552
box 22496 18552 22564 18752
use cut_M3M4_1x2 
transform 1 0 3644 0 1 18506
box 3644 18506 3712 18706
use cut_M2M3_1x2 
transform 1 0 12768 0 1 18506
box 12768 18506 12836 18706
use cut_M3M4_1x2 
transform 1 0 4484 0 1 18684
box 4484 18684 4552 18884
use cut_M2M3_1x2 
transform 1 0 12456 0 1 18684
box 12456 18684 12524 18884
use cut_M3M4_1x2 
transform 1 0 8284 0 1 18862
box 8284 18862 8352 19062
use cut_M2M3_1x2 
transform 1 0 12144 0 1 18862
box 12144 18862 12212 19062
use cut_M3M4_1x2 
transform 1 0 -156 0 1 19040
box -156 19040 -88 19240
use cut_M2M3_1x2 
transform 1 0 13080 0 1 19040
box 13080 19040 13148 19240
use cut_M3M4_1x2 
transform 1 0 12320 0 1 19218
box 12320 19218 12388 19418
use cut_M2M3_1x2 
transform 1 0 10508 0 1 19218
box 10508 19218 10576 19418
use cut_M3M4_1x2 
transform 1 0 16960 0 1 19396
box 16960 19396 17028 19596
use cut_M2M3_1x2 
transform 1 0 10820 0 1 19396
box 10820 19396 10888 19596
use cut_M3M4_1x2 
transform 1 0 9860 0 1 19574
box 9860 19574 9928 19774
use cut_M2M3_1x2 
transform 1 0 10352 0 1 19574
box 10352 19574 10420 19774
use cut_M3M4_1x2 
transform 1 0 14500 0 1 19752
box 14500 19752 14568 19952
use cut_M2M3_1x2 
transform 1 0 10664 0 1 19752
box 10664 19752 10732 19952
use cut_M3M4_1x2 
transform 1 0 580 0 1 19930
box 580 19930 648 20130
use cut_M2M3_1x2 
transform 1 0 9104 0 1 19930
box 9104 19930 9172 20130
use cut_M3M4_1x2 
transform 1 0 5220 0 1 20108
box 5220 20108 5288 20308
use cut_M2M3_1x2 
transform 1 0 9728 0 1 20108
box 9728 20108 9796 20308
use cut_M3M4_1x2 
transform 1 0 3040 0 1 20286
box 3040 20286 3108 20486
use cut_M2M3_1x2 
transform 1 0 9416 0 1 20286
box 9416 20286 9484 20486
use cut_M3M4_1x2 
transform 1 0 7680 0 1 20464
box 7680 20464 7748 20664
use cut_M2M3_1x2 
transform 1 0 10040 0 1 20464
box 10040 20464 10108 20664
use cut_M3M4_1x2 
transform 1 0 716 0 1 20642
box 716 20642 784 20842
use cut_M2M3_1x2 
transform 1 0 9260 0 1 20642
box 9260 20642 9328 20842
use cut_M3M4_1x2 
transform 1 0 7544 0 1 20820
box 7544 20820 7612 21020
use cut_M2M3_1x2 
transform 1 0 10196 0 1 20820
box 10196 20820 10264 21020
use cut_M3M4_1x2 
transform 1 0 5356 0 1 20998
box 5356 20998 5424 21198
use cut_M2M3_1x2 
transform 1 0 9884 0 1 20998
box 9884 20998 9952 21198
use cut_M3M4_1x2 
transform 1 0 2904 0 1 21176
box 2904 21176 2972 21376
use cut_M2M3_1x2 
transform 1 0 9572 0 1 21176
box 9572 21176 9640 21376
use cut_M3M4_1x2 
transform 1 0 10132 0 1 21354
box 10132 21354 10200 21554
use cut_M2M3_1x2 
transform 1 0 11832 0 1 21354
box 11832 21354 11900 21554
use cut_M3M4_1x2 
transform 1 0 12048 0 1 21532
box 12048 21532 12116 21732
use cut_M2M3_1x2 
transform 1 0 11676 0 1 21532
box 11676 21532 11744 21732
use cut_M3M4_1x2 
transform 1 0 14772 0 1 21710
box 14772 21710 14840 21910
use cut_M2M3_1x2 
transform 1 0 11520 0 1 21710
box 11520 21710 11588 21910
use cut_M3M4_1x2 
transform 1 0 7408 0 1 21888
box 7408 21888 7476 22088
use cut_M2M3_1x2 
transform 1 0 11988 0 1 21888
box 11988 21888 12056 22088
use cut_M3M4_1x2 
transform 1 0 2768 0 1 22066
box 2768 22066 2836 22266
use cut_M2M3_1x2 
transform 1 0 12612 0 1 22066
box 12612 22066 12680 22266
use cut_M3M4_1x2 
transform 1 0 852 0 1 22244
box 852 22244 920 22444
use cut_M2M3_1x2 
transform 1 0 12924 0 1 22244
box 12924 22244 12992 22444
use cut_M3M4_1x2 
transform 1 0 16688 0 1 22422
box 16688 22422 16756 22622
use cut_M2M3_1x2 
transform 1 0 11364 0 1 22422
box 11364 22422 11432 22622
use cut_M3M4_1x2 
transform 1 0 5492 0 1 22600
box 5492 22600 5560 22800
use cut_M2M3_1x2 
transform 1 0 12300 0 1 22600
box 12300 22600 12368 22800
<< labels >>
flabel m3 s -152 19170 -92 28628 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 12324 19348 12384 28642 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 16964 19526 17024 28642 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 9864 19704 9924 28642 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 14504 19882 14564 28642 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 5224 20238 5284 28642 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 3044 20416 3104 28642 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 7684 20594 7744 28642 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel m3 s 10208 46 10408 114 0 FreeSans 400 0 0 0 SAR_IP
port 9 nsew
flabel m3 s 11848 46 12048 114 0 FreeSans 400 0 0 0 SAR_IN
port 10 nsew
flabel locali s 10208 2450 10448 2510 0 FreeSans 400 0 0 0 SARN
port 11 nsew
flabel locali s 10208 1170 10448 1230 0 FreeSans 400 0 0 0 SARP
port 12 nsew
flabel locali s 18768 34152 19008 34212 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 19144 28642 19212 28842 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
flabel m2 s -152 23828 48 23896 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s -192 32792 48 32852 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 9248 450 9488 510 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel m3 s 1568 27752 1768 27952 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel m3 s 8168 0 8368 4800 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel m3 s 8888 0 9088 4800 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
<< end >>
