* SUN_PLL_BUF

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SUN_PLL_BUF_lpe.spi
.include ../../../design/SUN_PLL_SKY130NM.spice
#else
.include ../../../design/SUN_PLL_SKY130NM.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
*.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12
#else
*.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD  AVSS  dc {AVDD}
VPWR PWRUP_1V8 AVSS dc {AVDD}
VI VI 0 pwl 0 {AVDD/2} 10n {AVDD/2} 1u {AVDD}

IB 0 IBPSR_1U dc 1u

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
x2 IBPSR_1U AVDD PWRUP_1V8 AVSS SUN_PLL_BIAS
XDUT AVDD VO VI VO IBPSR_1U AVSS SUN_PLL_BUF
xh2 AVDD CK VO PWRUP_1V8 AVSS SUN_PLL_ROSC

*R1 VO 0 10k

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
*.probe v(*)
#else
.probe v(AVDD)  v(VI) v(VO) v(IBPSR_1U) v(AVSS) v(XDUT.VGP)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

#ifdef Debug
tran 10p 200n 1p
write
quit
#else
tran 10p 1u 1p
write
quit
#endif

.endc

.end


