magic
tech sky130A
magscale 1 2
timestamp 1660244192
<< checkpaint >>
rect 0 0 200 76
<< m2 >>
rect 0 0 200 76
<< m3 >>
rect 0 0 200 76
<< v2 >>
rect 12 6 188 70
<< labels >>
<< end >>
