magic
tech sky130A
magscale 1 2
timestamp 1660117866
<< checkpaint >>
rect -672 -672 36280 7392
<< locali >>
rect 36040 -672 36280 7392
rect -672 -672 36280 -432
rect -672 7152 36280 7392
rect -672 -672 -432 7392
rect 36040 -672 36280 7392
rect 216 -672 432 -88
rect -54 3190 270 3410
<< m3 >>
rect 18620 -672 18836 40
rect 18728 -40 35560 36
rect 18728 920 35560 996
rect 18728 1880 35560 1956
rect 18728 2840 35560 2916
rect 18728 3800 35560 3876
rect 18728 4760 35560 4836
rect 18728 5720 35560 5796
rect 35560 -40 35636 5796
<< m1 >>
rect 540 3190 762 3250
rect 762 2680 2068 2740
rect 762 3640 2068 3700
rect 762 4600 2068 4660
rect 762 5560 2068 5620
rect 762 6520 2068 6580
rect 762 2680 822 6596
<< m2 >>
rect 108 3190 334 3266
rect 334 760 2068 836
rect 334 1720 2068 1796
rect 334 760 410 3266
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO_12k xa30
transform 1 0 0 0 1 440
box 0 440 1928 4580
use CAP_LPF xb10
transform -1 0 35608 0 1 0
box 35608 0 69288 960
use CAP_LPF xb20
transform -1 0 35608 0 1 960
box 35608 960 69288 1920
use CAP_LPF xb30
transform -1 0 35608 0 1 1920
box 35608 1920 69288 2880
use CAP_LPF xb31
transform -1 0 35608 0 1 2880
box 35608 2880 69288 3840
use CAP_LPF xb32
transform -1 0 35608 0 1 3840
box 35608 3840 69288 4800
use CAP_LPF xb33
transform -1 0 35608 0 1 4800
box 35608 4800 69288 5760
use CAP_LPF xb34
transform -1 0 35608 0 1 5760
box 35608 5760 69288 6720
use cut_M1M4_2x1 
transform 1 0 18628 0 1 -672
box 18628 -672 18828 -596
use cut_M1M2_2x1 
transform 1 0 378 0 1 3190
box 378 3190 562 3258
use cut_M2M4_2x1 
transform 1 0 1968 0 1 2680
box 1968 2680 2168 2756
use cut_M2M4_2x1 
transform 1 0 1968 0 1 3640
box 1968 3640 2168 3716
use cut_M2M4_2x1 
transform 1 0 1968 0 1 4600
box 1968 4600 2168 4676
use cut_M2M4_2x1 
transform 1 0 1968 0 1 5560
box 1968 5560 2168 5636
use cut_M2M4_2x1 
transform 1 0 1968 0 1 6520
box 1968 6520 2168 6596
use cut_M1M3_2x1 
transform 1 0 -54 0 1 3190
box -54 3190 146 3266
use cut_M3M4_2x1 
transform 1 0 1968 0 1 760
box 1968 760 2168 836
use cut_M3M4_2x1 
transform 1 0 1968 0 1 1720
box 1968 1720 2168 1796
<< labels >>
flabel locali s 36040 -672 36280 7392 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s -54 3190 270 3410 0 FreeSans 400 0 0 0 VLPF
port 1 nsew
<< end >>
