magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect -648 0 22872 36734
<< m3 >>
rect 8580 17384 22702 17444
rect 8580 17724 22702 17784
rect 20562 18056 20622 24704
rect 20790 18056 20850 31744
rect 4722 18124 4782 27900
rect 5438 18294 5498 27900
rect 8682 18464 8742 27900
rect 1478 18634 1538 27900
rect 12078 18804 12138 27922
rect 16038 18974 16098 27922
rect 10078 19144 10138 27922
rect 14038 19314 14098 27922
rect 2158 19484 2218 27922
rect 6118 19654 6178 27922
rect 4158 19824 4218 27922
rect 8118 19994 8178 27922
rect 2294 20164 2354 29202
rect 7982 20334 8042 29202
rect 6254 20504 6314 29202
rect 4022 20674 4082 29202
rect 10350 20844 10410 30482
rect 11806 21014 11866 30482
rect 14310 21184 14370 30482
rect 7846 21354 7906 30482
rect 3886 21524 3946 30482
rect 2430 21694 2490 30482
rect 15766 21864 15826 30482
rect 6390 22034 6450 30482
<< m2 >>
rect 13572 16934 13632 17452
rect 8580 16934 8640 17792
rect 4722 18064 12816 18124
rect 5438 18234 12504 18294
rect 8682 18404 12192 18464
rect 1478 18574 13128 18634
rect 10496 18744 12138 18804
rect 10808 18914 16098 18974
rect 10078 19084 10400 19144
rect 10652 19254 14098 19314
rect 2158 19424 9152 19484
rect 6118 19594 9776 19654
rect 4158 19764 9464 19824
rect 8118 19934 10088 19994
rect 2294 20104 9308 20164
rect 7982 20274 10244 20334
rect 6254 20444 9932 20504
rect 4022 20614 9620 20674
rect 10350 20784 11880 20844
rect 11664 20954 11866 21014
rect 11508 21124 14370 21184
rect 7846 21294 12036 21354
rect 3886 21464 12660 21524
rect 2430 21634 12972 21694
rect 11352 21804 15826 21864
rect 6390 21974 12348 22034
<< m4 >>
rect 20562 17724 20622 18056
rect 20790 17384 20850 18056
<< m1 >>
rect 12756 16874 12816 18064
rect 12444 16874 12504 18234
rect 12132 16874 12192 18404
rect 13068 16874 13128 18574
rect 10496 16874 10556 18744
rect 10808 16874 10868 18914
rect 10340 16874 10400 19084
rect 10652 16874 10712 19254
rect 9092 16874 9152 19424
rect 9716 16874 9776 19594
rect 9404 16874 9464 19764
rect 10028 16874 10088 19934
rect 9248 16874 9308 20104
rect 10184 16874 10244 20274
rect 9872 16874 9932 20444
rect 9560 16874 9620 20614
rect 11820 16874 11880 20784
rect 11664 16874 11724 20954
rect 11508 16874 11568 21124
rect 11976 16874 12036 21294
rect 12600 16874 12660 21464
rect 12912 16874 12972 21634
rect 11352 16874 11412 21804
rect 12288 16874 12348 21974
use SARBSSW_CV XB1
transform -1 0 11112 0 1 0
box 11112 0 22872 4800
use SARBSSW_CV XB2
transform 1 0 11112 0 1 0
box 11112 0 22872 4800
use CDAC8_CV XDAC1
transform -1 0 10988 0 1 4970
box 10988 4970 21860 16934
use CDAC8_CV XDAC2
transform 1 0 11232 0 1 4970
box 11232 4970 22104 16934
use SARDIGEX4_CV XA0
transform 1 0 1212 0 1 22654
box 1212 22654 3192 35774
use SARDIGEX4_CV XA1
transform -1 0 5172 0 1 22654
box 5172 22654 7152 35774
use SARDIGEX4_CV XA2
transform 1 0 5172 0 1 22654
box 5172 22654 7152 35774
use SARDIGEX4_CV XA3
transform -1 0 9132 0 1 22654
box 9132 22654 11112 35774
use SARDIGEX4_CV XA4
transform 1 0 9132 0 1 22654
box 9132 22654 11112 35774
use SARDIGEX4_CV XA5
transform -1 0 13092 0 1 22654
box 13092 22654 15072 35774
use SARDIGEX4_CV XA6
transform 1 0 13092 0 1 22654
box 13092 22654 15072 35774
use SARDIGEX4_CV XA7
transform -1 0 17052 0 1 22654
box 17052 22654 19032 35774
use SARDIGEX4_CV XA8
transform 1 0 17052 0 1 22654
box 17052 22654 19032 35774
use SARCMPX1_CV XA20
transform -1 0 21012 0 1 22654
box 21012 22654 22992 36734
use cut_M3M4_1x2 
transform 1 0 13572 0 1 16934
box 13572 16934 13640 17118
use cut_M3M4_2x1 
transform 1 0 13572 0 1 17384
box 13572 17384 13756 17452
use cut_M3M4_1x2 
transform 1 0 8580 0 1 16934
box 8580 16934 8648 17118
use cut_M3M4_2x1 
transform 1 0 8580 0 1 17724
box 8580 17724 8764 17792
use cut_M2M4_2x1 
transform 1 0 20562 0 1 24704
box 20562 24704 20746 24772
use cut_M4M5_2x1 
transform 1 0 20562 0 1 17724
box 20562 17724 20746 17792
use cut_M4M5_1x2 
transform 1 0 20562 0 1 18056
box 20562 18056 20630 18240
use cut_M3M4_2x1 
transform 1 0 20666 0 1 31744
box 20666 31744 20850 31812
use cut_M2M3_2x1 
transform 1 0 20562 0 1 31744
box 20562 31744 20746 31812
use cut_M4M5_2x1 
transform 1 0 20790 0 1 17384
box 20790 17384 20974 17452
use cut_M4M5_1x2 
transform 1 0 20790 0 1 18056
box 20790 18056 20858 18240
use cut_M3M4_1x2 
transform 1 0 4718 0 1 18002
box 4718 18002 4786 18186
use cut_M2M3_1x2 
transform 1 0 12752 0 1 18002
box 12752 18002 12820 18186
use cut_M3M4_1x2 
transform 1 0 5434 0 1 18172
box 5434 18172 5502 18356
use cut_M2M3_1x2 
transform 1 0 12440 0 1 18172
box 12440 18172 12508 18356
use cut_M3M4_1x2 
transform 1 0 8678 0 1 18342
box 8678 18342 8746 18526
use cut_M2M3_1x2 
transform 1 0 12128 0 1 18342
box 12128 18342 12196 18526
use cut_M3M4_1x2 
transform 1 0 1474 0 1 18512
box 1474 18512 1542 18696
use cut_M2M3_1x2 
transform 1 0 13064 0 1 18512
box 13064 18512 13132 18696
use cut_M3M4_1x2 
transform 1 0 12074 0 1 18682
box 12074 18682 12142 18866
use cut_M2M3_1x2 
transform 1 0 10492 0 1 18682
box 10492 18682 10560 18866
use cut_M3M4_1x2 
transform 1 0 16034 0 1 18852
box 16034 18852 16102 19036
use cut_M2M3_1x2 
transform 1 0 10804 0 1 18852
box 10804 18852 10872 19036
use cut_M3M4_1x2 
transform 1 0 10074 0 1 19022
box 10074 19022 10142 19206
use cut_M2M3_1x2 
transform 1 0 10336 0 1 19022
box 10336 19022 10404 19206
use cut_M3M4_1x2 
transform 1 0 14034 0 1 19192
box 14034 19192 14102 19376
use cut_M2M3_1x2 
transform 1 0 10648 0 1 19192
box 10648 19192 10716 19376
use cut_M3M4_1x2 
transform 1 0 2154 0 1 19362
box 2154 19362 2222 19546
use cut_M2M3_1x2 
transform 1 0 9088 0 1 19362
box 9088 19362 9156 19546
use cut_M3M4_1x2 
transform 1 0 6114 0 1 19532
box 6114 19532 6182 19716
use cut_M2M3_1x2 
transform 1 0 9712 0 1 19532
box 9712 19532 9780 19716
use cut_M3M4_1x2 
transform 1 0 4154 0 1 19702
box 4154 19702 4222 19886
use cut_M2M3_1x2 
transform 1 0 9400 0 1 19702
box 9400 19702 9468 19886
use cut_M3M4_1x2 
transform 1 0 8114 0 1 19872
box 8114 19872 8182 20056
use cut_M2M3_1x2 
transform 1 0 10024 0 1 19872
box 10024 19872 10092 20056
use cut_M3M4_1x2 
transform 1 0 2290 0 1 20042
box 2290 20042 2358 20226
use cut_M2M3_1x2 
transform 1 0 9244 0 1 20042
box 9244 20042 9312 20226
use cut_M3M4_1x2 
transform 1 0 7978 0 1 20212
box 7978 20212 8046 20396
use cut_M2M3_1x2 
transform 1 0 10180 0 1 20212
box 10180 20212 10248 20396
use cut_M3M4_1x2 
transform 1 0 6250 0 1 20382
box 6250 20382 6318 20566
use cut_M2M3_1x2 
transform 1 0 9868 0 1 20382
box 9868 20382 9936 20566
use cut_M3M4_1x2 
transform 1 0 4018 0 1 20552
box 4018 20552 4086 20736
use cut_M2M3_1x2 
transform 1 0 9556 0 1 20552
box 9556 20552 9624 20736
use cut_M3M4_1x2 
transform 1 0 10346 0 1 20722
box 10346 20722 10414 20906
use cut_M2M3_1x2 
transform 1 0 11816 0 1 20722
box 11816 20722 11884 20906
use cut_M3M4_1x2 
transform 1 0 11802 0 1 20892
box 11802 20892 11870 21076
use cut_M2M3_1x2 
transform 1 0 11660 0 1 20892
box 11660 20892 11728 21076
use cut_M3M4_1x2 
transform 1 0 14306 0 1 21062
box 14306 21062 14374 21246
use cut_M2M3_1x2 
transform 1 0 11504 0 1 21062
box 11504 21062 11572 21246
use cut_M3M4_1x2 
transform 1 0 7842 0 1 21232
box 7842 21232 7910 21416
use cut_M2M3_1x2 
transform 1 0 11972 0 1 21232
box 11972 21232 12040 21416
use cut_M3M4_1x2 
transform 1 0 3882 0 1 21402
box 3882 21402 3950 21586
use cut_M2M3_1x2 
transform 1 0 12596 0 1 21402
box 12596 21402 12664 21586
use cut_M3M4_1x2 
transform 1 0 2426 0 1 21572
box 2426 21572 2494 21756
use cut_M2M3_1x2 
transform 1 0 12908 0 1 21572
box 12908 21572 12976 21756
use cut_M3M4_1x2 
transform 1 0 15762 0 1 21742
box 15762 21742 15830 21926
use cut_M2M3_1x2 
transform 1 0 11348 0 1 21742
box 11348 21742 11416 21926
use cut_M3M4_1x2 
transform 1 0 6386 0 1 21912
box 6386 21912 6454 22096
use cut_M2M3_1x2 
transform 1 0 12284 0 1 21912
box 12284 21912 12352 22096
<< labels >>
flabel m3 s 1478 18634 1538 27900 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 12078 18804 12138 27922 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 16038 18974 16098 27922 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 10078 19144 10138 27922 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 14038 19314 14098 27922 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 6118 19654 6178 27922 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 4158 19824 4218 27922 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8118 19994 8178 27922 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel m3 s 10302 46 10486 114 0 FreeSans 400 0 0 0 SAR_IP
port 9 nsew
flabel m3 s 11738 46 11922 114 0 FreeSans 400 0 0 0 SAR_IN
port 10 nsew
flabel locali s 10302 2450 10482 2510 0 FreeSans 400 0 0 0 SARN
port 11 nsew
flabel locali s 10302 1170 10482 1230 0 FreeSans 400 0 0 0 SARP
port 12 nsew
flabel locali s 17682 33424 17862 33484 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 17998 27922 18066 28106 0 FreeSans 400 0 0 0 D<0>
port 14 nsew
flabel m2 s 1478 23100 1662 23168 0 FreeSans 400 0 0 0 EN
port 15 nsew
flabel locali s 1482 32064 1662 32124 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 9522 450 9702 510 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 17 nsew
flabel m3 s 2862 27024 3046 27208 0 FreeSans 400 0 0 0 VREF
port 18 nsew
flabel m3 s 8618 0 8802 4800 0 FreeSans 400 0 0 0 AVDD
port 19 nsew
flabel m3 s 9158 0 9342 4800 0 FreeSans 400 0 0 0 AVSS
port 20 nsew
<< end >>
