magic
tech sky130A
magscale 1 2
timestamp 1658775803
<< checkpaint >>
rect 0 0 10152 1056
<< m1 >>
rect 108 -44 10116 44
rect 10044 44 10116 132
rect 108 132 9972 220
rect 10044 132 10116 220
rect 108 220 180 308
rect 10044 220 10116 308
rect 108 308 180 396
rect 252 308 10116 396
rect 108 396 180 484
rect 10044 396 10116 484
rect 108 484 9972 572
rect 10044 484 10116 572
rect 108 572 180 660
rect 10044 572 10116 660
rect 108 660 180 748
rect 252 660 10116 748
rect 108 748 180 836
rect 108 836 10116 924
<< m2 >>
rect 108 -44 10116 44
rect 10044 44 10116 132
rect 108 132 9972 220
rect 10044 132 10116 220
rect 108 220 180 308
rect 10044 220 10116 308
rect 108 308 180 396
rect 252 308 10116 396
rect 108 396 180 484
rect 10044 396 10116 484
rect 108 484 9972 572
rect 10044 484 10116 572
rect 108 572 180 660
rect 10044 572 10116 660
rect 108 660 180 748
rect 252 660 10116 748
rect 108 748 180 836
rect 108 836 10116 924
<< locali >>
rect 108 -44 10116 44
rect 10044 44 10116 132
rect 108 132 9972 220
rect 10044 132 10116 220
rect 108 220 180 308
rect 10044 220 10116 308
rect 108 308 180 396
rect 252 308 10116 396
rect 108 396 180 484
rect 10044 396 10116 484
rect 108 484 9972 572
rect 10044 484 10116 572
rect 108 572 180 660
rect 10044 572 10116 660
rect 108 660 180 748
rect 252 660 10116 748
rect 108 748 180 836
rect 108 836 10116 924
<< v1 >>
rect 9756 -35 9828 -26
rect 9756 -26 9828 -17
rect 9756 -17 9828 -8
rect 9756 -8 9828 0
rect 9756 0 9828 8
rect 9756 8 9828 17
rect 9756 17 9828 26
rect 9756 26 9828 35
rect 9828 -35 9900 -26
rect 9828 -26 9900 -17
rect 9828 -17 9900 -8
rect 9828 -8 9900 0
rect 9828 0 9900 8
rect 9828 8 9900 17
rect 9828 17 9900 26
rect 9828 26 9900 35
rect 9900 -35 9972 -26
rect 9900 -26 9972 -17
rect 9900 -17 9972 -8
rect 9900 -8 9972 0
rect 9900 0 9972 8
rect 9900 8 9972 17
rect 9900 17 9972 26
rect 9900 26 9972 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 9756 316 9828 325
rect 9756 325 9828 334
rect 9756 334 9828 343
rect 9756 343 9828 352
rect 9756 352 9828 360
rect 9756 360 9828 369
rect 9756 369 9828 378
rect 9756 378 9828 387
rect 9828 316 9900 325
rect 9828 325 9900 334
rect 9828 334 9900 343
rect 9828 343 9900 352
rect 9828 352 9900 360
rect 9828 360 9900 369
rect 9828 369 9900 378
rect 9828 378 9900 387
rect 9900 316 9972 325
rect 9900 325 9972 334
rect 9900 334 9972 343
rect 9900 343 9972 352
rect 9900 352 9972 360
rect 9900 360 9972 369
rect 9900 369 9972 378
rect 9900 378 9972 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 9756 668 9828 677
rect 9756 677 9828 686
rect 9756 686 9828 695
rect 9756 695 9828 704
rect 9756 704 9828 712
rect 9756 712 9828 721
rect 9756 721 9828 730
rect 9756 730 9828 739
rect 9828 668 9900 677
rect 9828 677 9900 686
rect 9828 686 9900 695
rect 9828 695 9900 704
rect 9828 704 9900 712
rect 9828 712 9900 721
rect 9828 721 9900 730
rect 9828 730 9900 739
rect 9900 668 9972 677
rect 9900 677 9972 686
rect 9900 686 9972 695
rect 9900 695 9972 704
rect 9900 704 9972 712
rect 9900 712 9972 721
rect 9900 721 9972 730
rect 9900 730 9972 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 9756 -35 9828 -26
rect 9756 -26 9828 -17
rect 9756 -17 9828 -8
rect 9756 -8 9828 0
rect 9756 0 9828 8
rect 9756 8 9828 17
rect 9756 17 9828 26
rect 9756 26 9828 35
rect 9828 -35 9900 -26
rect 9828 -26 9900 -17
rect 9828 -17 9900 -8
rect 9828 -8 9900 0
rect 9828 0 9900 8
rect 9828 8 9900 17
rect 9828 17 9900 26
rect 9828 26 9900 35
rect 9900 -35 9972 -26
rect 9900 -26 9972 -17
rect 9900 -17 9972 -8
rect 9900 -8 9972 0
rect 9900 0 9972 8
rect 9900 8 9972 17
rect 9900 17 9972 26
rect 9900 26 9972 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 9756 316 9828 325
rect 9756 325 9828 334
rect 9756 334 9828 343
rect 9756 343 9828 352
rect 9756 352 9828 360
rect 9756 360 9828 369
rect 9756 369 9828 378
rect 9756 378 9828 387
rect 9828 316 9900 325
rect 9828 325 9900 334
rect 9828 334 9900 343
rect 9828 343 9900 352
rect 9828 352 9900 360
rect 9828 360 9900 369
rect 9828 369 9900 378
rect 9828 378 9900 387
rect 9900 316 9972 325
rect 9900 325 9972 334
rect 9900 334 9972 343
rect 9900 343 9972 352
rect 9900 352 9972 360
rect 9900 360 9972 369
rect 9900 369 9972 378
rect 9900 378 9972 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 9756 668 9828 677
rect 9756 677 9828 686
rect 9756 686 9828 695
rect 9756 695 9828 704
rect 9756 704 9828 712
rect 9756 712 9828 721
rect 9756 721 9828 730
rect 9756 730 9828 739
rect 9828 668 9900 677
rect 9828 677 9900 686
rect 9828 686 9900 695
rect 9828 695 9900 704
rect 9828 704 9900 712
rect 9828 712 9900 721
rect 9828 721 9900 730
rect 9828 730 9900 739
rect 9900 668 9972 677
rect 9900 677 9972 686
rect 9900 686 9972 695
rect 9900 695 9972 704
rect 9900 704 9972 712
rect 9900 712 9972 721
rect 9900 721 9972 730
rect 9900 730 9972 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 9756 -35 9828 -26
rect 9756 -26 9828 -17
rect 9756 -17 9828 -8
rect 9756 -8 9828 0
rect 9756 0 9828 8
rect 9756 8 9828 17
rect 9756 17 9828 26
rect 9756 26 9828 35
rect 9828 -35 9900 -26
rect 9828 -26 9900 -17
rect 9828 -17 9900 -8
rect 9828 -8 9900 0
rect 9828 0 9900 8
rect 9828 8 9900 17
rect 9828 17 9900 26
rect 9828 26 9900 35
rect 9900 -35 9972 -26
rect 9900 -26 9972 -17
rect 9900 -17 9972 -8
rect 9900 -8 9972 0
rect 9900 0 9972 8
rect 9900 8 9972 17
rect 9900 17 9972 26
rect 9900 26 9972 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 9756 316 9828 325
rect 9756 325 9828 334
rect 9756 334 9828 343
rect 9756 343 9828 352
rect 9756 352 9828 360
rect 9756 360 9828 369
rect 9756 369 9828 378
rect 9756 378 9828 387
rect 9828 316 9900 325
rect 9828 325 9900 334
rect 9828 334 9900 343
rect 9828 343 9900 352
rect 9828 352 9900 360
rect 9828 360 9900 369
rect 9828 369 9900 378
rect 9828 378 9900 387
rect 9900 316 9972 325
rect 9900 325 9972 334
rect 9900 334 9972 343
rect 9900 343 9972 352
rect 9900 352 9972 360
rect 9900 360 9972 369
rect 9900 369 9972 378
rect 9900 378 9972 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 9756 668 9828 677
rect 9756 677 9828 686
rect 9756 686 9828 695
rect 9756 695 9828 704
rect 9756 704 9828 712
rect 9756 712 9828 721
rect 9756 721 9828 730
rect 9756 730 9828 739
rect 9828 668 9900 677
rect 9828 677 9900 686
rect 9828 686 9900 695
rect 9828 695 9900 704
rect 9828 704 9900 712
rect 9828 712 9900 721
rect 9828 721 9900 730
rect 9828 730 9900 739
rect 9900 668 9972 677
rect 9900 677 9972 686
rect 9900 686 9972 695
rect 9900 695 9972 704
rect 9900 704 9972 712
rect 9900 712 9972 721
rect 9900 721 9972 730
rect 9900 730 9972 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 10116 44
rect 108 -44 10116 44
rect 10044 44 10116 132
rect 108 132 9756 220
rect 9828 132 9972 220
rect 10044 132 10116 220
rect 108 220 180 308
rect 10044 220 10116 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 10116 396
rect 108 396 180 484
rect 10044 396 10116 484
rect 108 484 9972 572
rect 10044 484 10116 572
rect 108 572 180 660
rect 10044 572 10116 660
rect 108 660 180 748
rect 252 660 10116 748
rect 108 748 180 836
rect 108 836 10116 924
rect 108 836 10116 924
<< rm3 >>
rect 9756 132 9828 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 10116 44 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel m3 s 108 836 10116 924 0 FreeSans 400 0 0 0 A
port 1 nsew
<< end >>
