magic
tech sky130A
magscale 1 2
timestamp 1659197050
<< checkpaint >>
rect 0 -1788 30240 8336
<< locali >>
rect 0 -720 30240 -520
rect 0 -720 30240 -520
rect 0 -1440 30240 -1240
rect 0 -1440 30240 -1240
rect 0 -1788 30240 -1728
rect 0 -1788 30240 -1728
rect 0 6480 30240 6540
rect 0 6480 30240 6540
rect 0 6684 30240 6744
rect 0 6684 30240 6744
rect 0 6816 956 6876
rect 0 6816 956 6876
rect 0 6948 4268 7008
rect 0 6948 4268 7008
rect 0 7080 5996 7140
rect 0 7080 5996 7140
rect 0 7212 9308 7272
rect 0 7212 9308 7272
rect 0 7344 11036 7404
rect 0 7344 11036 7404
rect 0 7476 14348 7536
rect 0 7476 14348 7536
rect 0 7608 16076 7668
rect 0 7608 16076 7668
rect 0 7740 19388 7800
rect 0 7740 19388 7800
rect 0 7872 21116 7932
rect 0 7872 21116 7932
rect 0 8004 24428 8064
rect 0 8004 24428 8064
rect 0 8136 26156 8196
rect 0 8136 26156 8196
rect 0 8268 29468 8328
rect 0 8268 29468 8328
rect 324 1906 540 1966
rect 4500 1906 4716 1966
rect 5364 1906 5580 1966
rect 9540 1906 9756 1966
rect 10404 1906 10620 1966
rect 14580 1906 14796 1966
rect 15444 1906 15660 1966
rect 19620 1906 19836 1966
rect 20484 1906 20700 1966
rect 24660 1906 24876 1966
rect 25524 1906 25740 1966
rect 29700 1906 29916 1966
<< m3 >>
rect 756 -720 956 6336
rect 4084 -720 4284 6336
rect 5796 -720 5996 6336
rect 9124 -720 9324 6336
rect 10836 -720 11036 6336
rect 14164 -720 14364 6336
rect 15876 -720 16076 6336
rect 19204 -720 19404 6336
rect 20916 -720 21116 6336
rect 24244 -720 24444 6336
rect 25956 -720 26156 6336
rect 29284 -720 29484 6336
rect 1548 -1440 1748 6336
rect 3292 -1440 3492 6336
rect 6588 -1440 6788 6336
rect 8332 -1440 8532 6336
rect 11628 -1440 11828 6336
rect 13372 -1440 13572 6336
rect 16668 -1440 16868 6336
rect 18412 -1440 18612 6336
rect 21708 -1440 21908 6336
rect 23452 -1440 23652 6336
rect 26748 -1440 26948 6336
rect 28492 -1440 28692 6336
<< m1 >>
rect 402 -1788 462 910
rect 4578 -1788 4638 910
rect 5442 -1788 5502 910
rect 9618 -1788 9678 910
rect 10482 -1788 10542 910
rect 14658 -1788 14718 910
rect 15522 -1788 15582 910
rect 19698 -1788 19758 910
rect 20562 -1788 20622 910
rect 24738 -1788 24798 910
rect 25602 -1788 25662 910
rect 29778 -1788 29838 910
rect 402 6130 462 6540
rect 4578 6130 4638 6540
rect 5442 6130 5502 6540
rect 9618 6130 9678 6540
rect 10482 6130 10542 6540
rect 14658 6130 14718 6540
rect 15522 6130 15582 6540
rect 19698 6130 19758 6540
rect 20562 6130 20622 6540
rect 24738 6130 24798 6540
rect 25602 6130 25662 6540
rect 29778 6130 29838 6540
rect 2058 6130 2118 6744
rect 2922 6130 2982 6744
rect 7098 6130 7158 6744
rect 7962 6130 8022 6744
rect 12138 6130 12198 6744
rect 13002 6130 13062 6744
rect 17178 6130 17238 6744
rect 18042 6130 18102 6744
rect 22218 6130 22278 6744
rect 23082 6130 23142 6744
rect 27258 6130 27318 6744
rect 28122 6130 28182 6744
rect 834 6218 894 6876
rect 4146 6218 4206 7008
rect 5874 6218 5934 7140
rect 9186 6218 9246 7272
rect 10914 6218 10974 7404
rect 14226 6218 14286 7536
rect 15954 6218 16014 7668
rect 19266 6218 19326 7800
rect 20994 6218 21054 7932
rect 24306 6218 24366 8064
rect 26034 6218 26094 8196
rect 29346 6218 29406 8328
use SUNTR_DFTRIX1_CV XA0
transform 1 0 0 0 1 0
box 0 0 2520 6336
use SUNTR_DFTRIX1_CV XB1
transform -1 0 5040 0 1 0
box 5040 0 7560 6336
use SUNTR_DFTRIX1_CV XC2
transform 1 0 5040 0 1 0
box 5040 0 7560 6336
use SUNTR_DFTRIX1_CV XD3
transform -1 0 10080 0 1 0
box 10080 0 12600 6336
use SUNTR_DFTRIX1_CV XE4
transform 1 0 10080 0 1 0
box 10080 0 12600 6336
use SUNTR_DFTRIX1_CV XF5
transform -1 0 15120 0 1 0
box 15120 0 17640 6336
use SUNTR_DFTRIX1_CV XG6
transform 1 0 15120 0 1 0
box 15120 0 17640 6336
use SUNTR_DFTRIX1_CV XH7
transform -1 0 20160 0 1 0
box 20160 0 22680 6336
use SUNTR_DFTRIX1_CV XI8
transform 1 0 20160 0 1 0
box 20160 0 22680 6336
use SUNTR_DFTRIX1_CV XJ9
transform -1 0 25200 0 1 0
box 25200 0 27720 6336
use SUNTR_DFTRIX1_CV XK10
transform 1 0 25200 0 1 0
box 25200 0 27720 6336
use SUNTR_DFTRIX1_CV XL11
transform -1 0 30240 0 1 0
box 30240 0 32760 6336
use SUNTR_cut_M1M4_2x2 
transform 1 0 756 0 1 -720
box 756 -720 956 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 4084 0 1 -720
box 4084 -720 4284 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 5796 0 1 -720
box 5796 -720 5996 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 9124 0 1 -720
box 9124 -720 9324 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 10836 0 1 -720
box 10836 -720 11036 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 14164 0 1 -720
box 14164 -720 14364 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 15876 0 1 -720
box 15876 -720 16076 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 19204 0 1 -720
box 19204 -720 19404 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 20916 0 1 -720
box 20916 -720 21116 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 24244 0 1 -720
box 24244 -720 24444 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 25956 0 1 -720
box 25956 -720 26156 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 29284 0 1 -720
box 29284 -720 29484 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 1548 0 1 -1440
box 1548 -1440 1748 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 3292 0 1 -1440
box 3292 -1440 3492 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 6588 0 1 -1440
box 6588 -1440 6788 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 8332 0 1 -1440
box 8332 -1440 8532 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 11628 0 1 -1440
box 11628 -1440 11828 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 13372 0 1 -1440
box 13372 -1440 13572 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 16668 0 1 -1440
box 16668 -1440 16868 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 18412 0 1 -1440
box 18412 -1440 18612 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 21708 0 1 -1440
box 21708 -1440 21908 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 23452 0 1 -1440
box 23452 -1440 23652 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 26748 0 1 -1440
box 26748 -1440 26948 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 28492 0 1 -1440
box 28492 -1440 28692 -1240
use SUNTR_cut_M1M2_2x1 
transform 1 0 340 0 1 850
box 340 850 524 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 340 0 1 -1788
box 340 -1788 524 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 4516 0 1 850
box 4516 850 4700 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 4516 0 1 -1788
box 4516 -1788 4700 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 5380 0 1 850
box 5380 850 5564 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 5380 0 1 -1788
box 5380 -1788 5564 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 9556 0 1 850
box 9556 850 9740 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 9556 0 1 -1788
box 9556 -1788 9740 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 10420 0 1 850
box 10420 850 10604 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 10420 0 1 -1788
box 10420 -1788 10604 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 14596 0 1 850
box 14596 850 14780 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 14596 0 1 -1788
box 14596 -1788 14780 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 15460 0 1 850
box 15460 850 15644 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 15460 0 1 -1788
box 15460 -1788 15644 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 19636 0 1 850
box 19636 850 19820 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 19636 0 1 -1788
box 19636 -1788 19820 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 20500 0 1 850
box 20500 850 20684 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 20500 0 1 -1788
box 20500 -1788 20684 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 24676 0 1 850
box 24676 850 24860 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 24676 0 1 -1788
box 24676 -1788 24860 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 25540 0 1 850
box 25540 850 25724 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 25540 0 1 -1788
box 25540 -1788 25724 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 29716 0 1 850
box 29716 850 29900 918
use SUNTR_cut_M1M2_2x1 
transform 1 0 29716 0 1 -1788
box 29716 -1788 29900 -1720
use SUNTR_cut_M1M2_2x1 
transform 1 0 340 0 1 6130
box 340 6130 524 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 340 0 1 6480
box 340 6480 524 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 4516 0 1 6130
box 4516 6130 4700 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 4516 0 1 6480
box 4516 6480 4700 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 5380 0 1 6130
box 5380 6130 5564 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 5380 0 1 6480
box 5380 6480 5564 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 9556 0 1 6130
box 9556 6130 9740 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 9556 0 1 6480
box 9556 6480 9740 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 10420 0 1 6130
box 10420 6130 10604 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 10420 0 1 6480
box 10420 6480 10604 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 14596 0 1 6130
box 14596 6130 14780 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 14596 0 1 6480
box 14596 6480 14780 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 15460 0 1 6130
box 15460 6130 15644 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 15460 0 1 6480
box 15460 6480 15644 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 19636 0 1 6130
box 19636 6130 19820 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 19636 0 1 6480
box 19636 6480 19820 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 20500 0 1 6130
box 20500 6130 20684 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 20500 0 1 6480
box 20500 6480 20684 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 24676 0 1 6130
box 24676 6130 24860 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 24676 0 1 6480
box 24676 6480 24860 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 25540 0 1 6130
box 25540 6130 25724 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 25540 0 1 6480
box 25540 6480 25724 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 29716 0 1 6130
box 29716 6130 29900 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 29716 0 1 6480
box 29716 6480 29900 6548
use SUNTR_cut_M1M2_2x1 
transform 1 0 1996 0 1 6130
box 1996 6130 2180 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 1996 0 1 6684
box 1996 6684 2180 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 2860 0 1 6130
box 2860 6130 3044 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 2860 0 1 6684
box 2860 6684 3044 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 7036 0 1 6130
box 7036 6130 7220 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 7036 0 1 6684
box 7036 6684 7220 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 7900 0 1 6130
box 7900 6130 8084 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 7900 0 1 6684
box 7900 6684 8084 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 12076 0 1 6130
box 12076 6130 12260 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 12076 0 1 6684
box 12076 6684 12260 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 12940 0 1 6130
box 12940 6130 13124 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 12940 0 1 6684
box 12940 6684 13124 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 17116 0 1 6130
box 17116 6130 17300 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 17116 0 1 6684
box 17116 6684 17300 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 17980 0 1 6130
box 17980 6130 18164 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 17980 0 1 6684
box 17980 6684 18164 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 22156 0 1 6130
box 22156 6130 22340 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 22156 0 1 6684
box 22156 6684 22340 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 23020 0 1 6130
box 23020 6130 23204 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 23020 0 1 6684
box 23020 6684 23204 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 27196 0 1 6130
box 27196 6130 27380 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 27196 0 1 6684
box 27196 6684 27380 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 28060 0 1 6130
box 28060 6130 28244 6198
use SUNTR_cut_M1M2_2x1 
transform 1 0 28060 0 1 6684
box 28060 6684 28244 6752
use SUNTR_cut_M1M2_2x1 
transform 1 0 772 0 1 6218
box 772 6218 956 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 772 0 1 6816
box 772 6816 956 6884
use SUNTR_cut_M1M2_2x1 
transform 1 0 4084 0 1 6218
box 4084 6218 4268 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 4084 0 1 6948
box 4084 6948 4268 7016
use SUNTR_cut_M1M2_2x1 
transform 1 0 5812 0 1 6218
box 5812 6218 5996 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 5812 0 1 7080
box 5812 7080 5996 7148
use SUNTR_cut_M1M2_2x1 
transform 1 0 9124 0 1 6218
box 9124 6218 9308 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 9124 0 1 7212
box 9124 7212 9308 7280
use SUNTR_cut_M1M2_2x1 
transform 1 0 10852 0 1 6218
box 10852 6218 11036 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 10852 0 1 7344
box 10852 7344 11036 7412
use SUNTR_cut_M1M2_2x1 
transform 1 0 14164 0 1 6218
box 14164 6218 14348 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 14164 0 1 7476
box 14164 7476 14348 7544
use SUNTR_cut_M1M2_2x1 
transform 1 0 15892 0 1 6218
box 15892 6218 16076 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 15892 0 1 7608
box 15892 7608 16076 7676
use SUNTR_cut_M1M2_2x1 
transform 1 0 19204 0 1 6218
box 19204 6218 19388 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 19204 0 1 7740
box 19204 7740 19388 7808
use SUNTR_cut_M1M2_2x1 
transform 1 0 20932 0 1 6218
box 20932 6218 21116 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 20932 0 1 7872
box 20932 7872 21116 7940
use SUNTR_cut_M1M2_2x1 
transform 1 0 24244 0 1 6218
box 24244 6218 24428 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 24244 0 1 8004
box 24244 8004 24428 8072
use SUNTR_cut_M1M2_2x1 
transform 1 0 25972 0 1 6218
box 25972 6218 26156 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 25972 0 1 8136
box 25972 8136 26156 8204
use SUNTR_cut_M1M2_2x1 
transform 1 0 29284 0 1 6218
box 29284 6218 29468 6286
use SUNTR_cut_M1M2_2x1 
transform 1 0 29284 0 1 8268
box 29284 8268 29468 8336
<< labels >>
flabel locali s 0 -720 30240 -520 0 FreeSans 400 0 0 0 AVSS
port 29 nsew
flabel locali s 0 -1440 30240 -1240 0 FreeSans 400 0 0 0 AVDD
port 28 nsew
flabel locali s 0 -1788 30240 -1728 0 FreeSans 400 0 0 0 CK
port 13 nsew
flabel locali s 0 6480 30240 6540 0 FreeSans 400 0 0 0 C
port 14 nsew
flabel locali s 0 6684 30240 6744 0 FreeSans 400 0 0 0 CN
port 15 nsew
flabel locali s 0 6816 956 6876 0 FreeSans 400 0 0 0 Y<11>
port 16 nsew
flabel locali s 0 6948 4268 7008 0 FreeSans 400 0 0 0 Y<10>
port 17 nsew
flabel locali s 0 7080 5996 7140 0 FreeSans 400 0 0 0 Y<9>
port 18 nsew
flabel locali s 0 7212 9308 7272 0 FreeSans 400 0 0 0 Y<8>
port 19 nsew
flabel locali s 0 7344 11036 7404 0 FreeSans 400 0 0 0 Y<7>
port 20 nsew
flabel locali s 0 7476 14348 7536 0 FreeSans 400 0 0 0 Y<6>
port 21 nsew
flabel locali s 0 7608 16076 7668 0 FreeSans 400 0 0 0 Y<5>
port 22 nsew
flabel locali s 0 7740 19388 7800 0 FreeSans 400 0 0 0 Y<4>
port 23 nsew
flabel locali s 0 7872 21116 7932 0 FreeSans 400 0 0 0 Y<3>
port 24 nsew
flabel locali s 0 8004 24428 8064 0 FreeSans 400 0 0 0 Y<2>
port 25 nsew
flabel locali s 0 8136 26156 8196 0 FreeSans 400 0 0 0 Y<1>
port 26 nsew
flabel locali s 0 8268 29468 8328 0 FreeSans 400 0 0 0 Y<0>
port 27 nsew
flabel locali s 324 1906 540 1966 0 FreeSans 400 0 0 0 D<11>
port 1 nsew
flabel locali s 4500 1906 4716 1966 0 FreeSans 400 0 0 0 D<10>
port 2 nsew
flabel locali s 5364 1906 5580 1966 0 FreeSans 400 0 0 0 D<9>
port 3 nsew
flabel locali s 9540 1906 9756 1966 0 FreeSans 400 0 0 0 D<8>
port 4 nsew
flabel locali s 10404 1906 10620 1966 0 FreeSans 400 0 0 0 D<7>
port 5 nsew
flabel locali s 14580 1906 14796 1966 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel locali s 15444 1906 15660 1966 0 FreeSans 400 0 0 0 D<5>
port 7 nsew
flabel locali s 19620 1906 19836 1966 0 FreeSans 400 0 0 0 D<4>
port 8 nsew
flabel locali s 20484 1906 20700 1966 0 FreeSans 400 0 0 0 D<3>
port 9 nsew
flabel locali s 24660 1906 24876 1966 0 FreeSans 400 0 0 0 D<2>
port 10 nsew
flabel locali s 25524 1906 25740 1966 0 FreeSans 400 0 0 0 D<1>
port 11 nsew
flabel locali s 29700 1906 29916 1966 0 FreeSans 400 0 0 0 D<0>
port 12 nsew
<< end >>
