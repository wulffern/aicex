* Transistor library

.SUBCKT PCHL D G S B
XM1 D G S B sky130_fd_pr__pfet_01v8_lvt  w=0.88  l=0.18
.ENDS

.SUBCKT NCHL D G S B
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt  w=0.88  l=0.18
.ENDS

.SUBCKT NCHCM D G S B
XM0 N0 G S B NCHL
XM1 N1 G N0 B NCHL
XM4 N2 G N1 B NCHL
XM5 D G N2 B NCHL
.ENDS

.SUBCKT PCHCM D G S B
XM0 N0 G S B PCHL
XM1 N1 G N0 B PCHL
XM4 N2 G N1 B PCHL
XM5 D G N2 B PCHL
.ENDS

.SUBCKT NCHA D G S B
XM0 D G S B NCHL
XM1 S G D B NCHL
.ENDS

.SUBCKT PCHA D G S B
XM0 D G S B PCHL
XM1 S G D B PCHL
.ENDS

.SUBCKT NCHCM2 D G S B
XM0 D G S B NCHCM
XM1 S G D B NCHCM
.ENDS

.SUBCKT PCHCM2 D G S B
XM0 D G S B PCHCM
XM1 S G D B PCHCM
.ENDS


.SUBCKT TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS NCHL
XMP1 AVDD AVDD AVDD AVDD PCHL
.ENDS

.SUBCKT TIEH_CV Y AVDD AVSS
XMN0 A A AVSS AVSS NCHL
XMP0 Y A AVDD AVDD PCHL
.ENDS

.SUBCKT TIEL_CV Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMP0 A A AVDD AVDD PCHL
.ENDS

.SUBCKT IVX1_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMP0 Y A AVDD AVDD PCHL
.ENDS

.SUBCKT IVX2_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMN1 AVSS A Y AVSS NCHL
XMP0 Y A AVDD AVDD PCHL
XMP1 AVDD A Y AVDD PCHL
.ENDS

.SUBCKT IVX4_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMN1 AVSS A Y AVSS NCHL
XMN2 Y A AVSS AVSS NCHL
XMN3 AVSS A Y AVSS NCHL
XMP0 Y A AVDD AVDD PCHL
XMP1 AVDD A Y AVDD PCHL
XMP2 Y A AVDD AVDD PCHL
XMP3 AVDD A Y AVDD PCHL
.ENDS

.SUBCKT IVX8_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMN1 AVSS A Y AVSS NCHL
XMN2 Y A AVSS AVSS NCHL
XMN3 AVSS A Y AVSS NCHL
XMN4 Y A AVSS AVSS NCHL
XMN5 AVSS A Y AVSS NCHL
XMN6 Y A AVSS AVSS NCHL
XMN7 AVSS A Y AVSS NCHL
XMP0 Y A AVDD AVDD PCHL
XMP1 AVDD A Y AVDD PCHL
XMP2 Y A AVDD AVDD PCHL
XMP3 AVDD A Y AVDD PCHL
XMP4 Y A AVDD AVDD PCHL
XMP5 AVDD A Y AVDD PCHL
XMP6 Y A AVDD AVDD PCHL
XMP7 AVDD A Y AVDD PCHL
.ENDS

.SUBCKT BFX1_CV A Y AVDD AVSS
XMN0 AVSS A B AVSS NCHL
XMN1 Y B AVSS AVSS NCHL
XMP0 AVDD A B AVDD PCHL
XMP1 Y B AVDD AVDD PCHL
.ENDS

.SUBCKT NRX1_CV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMN1 AVSS B Y AVSS NCHL
XMP0 N1 A AVDD AVDD PCHL
XMP1 Y B N1 AVDD PCHL
.ENDS

.SUBCKT NDX1_CV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS NCHL
XMN1 Y B N1 AVSS NCHL
XMP0 Y A AVDD AVDD PCHL
XMP1 AVDD B Y AVDD PCHL
.ENDS

.SUBCKT ORX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ORX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ORX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NRX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT ANX8_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS NDX1_CV
XA2 YN Y AVDD AVSS IVX1_CV
.ENDS

.SUBCKT IVTRIX1_CV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS NCHL
XMN1 Y C N1 AVSS NCHL
XMP0 N2 A AVDD AVDD PCHL
XMP1 Y CN N2 AVDD PCHL
.ENDS

.SUBCKT NDTRIX1_CV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS NCHL
XMN0 N2 A N1 AVSS NCHL
XMN1 Y C N2 AVSS NCHL
XMP2 AVDD RN N2 AVDD PCHL
XMP0 N2 A AVDD AVDD PCHL
XMP1 Y CN N2 AVDD PCHL
.ENDS

.SUBCKT DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS IVTRIX1_CV
XA5 A0 A1 AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS NDTRIX1_CV
XA8 QN Q AVDD AVSS IVX1_CV
.ENDS


.SUBCKT DFSRQNX1_CV D CK S R Q QN AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA0a R RN AVDD AVSS IVX1_CV
XA1 CK RN CKN AVDD AVSS NDX1_CV
XA2 CKN CKB AVDD AVSS IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS IVTRIX1_CV
XA5 A0 A1 AVDD AVSS IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS NDTRIX1_CV
XA8 QN Q AVDD AVSS IVX1_CV
.ENDS



.SUBCKT SCX1_CV A Y AVDD AVSS
XA2 N1 A AVSS AVSS NCHL
XA3 SCO A N1 AVSS NCHL
XA4a AVDD SCO N1 AVSS NCHL
XA4b AVDD SCO N1 AVSS NCHL
XA5 Y SCO AVSS AVSS NCHL
XB0 N2 A AVDD AVDD PCHL
XB1 SCO A N2 AVDD PCHL
XB3a N2 SCO AVSS AVDD PCHL
XB3b N2 SCO AVSS AVDD PCHL
XB4 Y SCO AVDD AVDD PCHL
.ENDS

.SUBCKT SWX2_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMN1 AVSS A Y AVSS NCHL
XMP0 Y A VREF AVDD PCHL
XMP1 VREF A Y AVDD PCHL
.ENDS

.SUBCKT SWX4_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS NCHL
XMN1 AVSS A Y AVSS NCHL
XMN2 Y A AVSS AVSS NCHL
XMN3 AVSS A Y AVSS NCHL
XMP0 Y A VREF AVDD PCHL
XMP1 VREF A Y AVDD PCHL
XMP2 Y A VREF AVDD PCHL
XMP3 VREF A Y AVDD PCHL
.ENDS

.SUBCKT TGPD_CV C A B AVDD AVSS
XMN0 AVSS C CN AVSS NCHL
XMN1 B C AVSS AVSS NCHL
XMN2 A CN B AVSS NCHL
XMP0 AVDD C CN AVDD PCHL
XMP1_DMY B AVDD AVDD AVDD PCHL
XMP2 A C B AVDD PCHL
.ENDS

.SUBCKT SUN_TR AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 Y1 AVDD AVSS TIEH_CV
XA2 Y2 AVDD AVSS TIEL_CV
XB0 AVDD AVSS TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS IVX1_CV
XB4 A4 Y4 AVDD AVSS IVX2_CV
XB5 A5 Y5 AVDD AVSS IVX4_CV
XB6 A6 Y6 AVDD AVSS IVX8_CV
XC0 AVDD AVSS TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS BFX1_CV
XD0 AVDD AVSS TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS ANX1_CV
XE0 AVDD AVSS TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SCX1_CV
XF0 AVDD AVSS TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS TGPD_CV
.ENDS

