magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 116 0 10988 11964
<< m1 >>
rect 1836 4596 1896 11904
rect 1680 132 1740 11904
rect 1524 9060 1584 11904
rect 1368 1620 1428 11904
rect 1212 3328 1272 11904
rect 1056 7792 1116 11904
rect 900 7572 960 11904
rect 744 8232 804 11904
rect 588 3768 648 11904
rect 432 3988 492 11904
rect 276 3548 336 11904
rect 120 4208 180 11904
<< m2 >>
rect 2028 4654 1896 4722
rect 2028 5754 1896 5822
rect 2028 5094 1896 5162
rect 2028 5534 1896 5602
rect 2028 5314 1896 5382
rect 2028 4874 1896 4942
rect 2028 4654 1896 4722
rect 2028 5754 1896 5822
rect 2028 5094 1896 5162
rect 2028 5534 1896 5602
rect 2028 5314 1896 5382
rect 2028 4874 1896 4942
rect 2028 4654 1896 4722
rect 2028 5754 1896 5822
rect 2028 5094 1896 5162
rect 2028 5534 1896 5602
rect 2028 5314 1896 5382
rect 2028 4874 1896 4942
rect 2028 4654 1896 4722
rect 2028 5754 1896 5822
rect 2028 5094 1896 5162
rect 2028 5534 1896 5602
rect 2028 5314 1896 5382
rect 2028 4874 1896 4942
rect 2028 4654 1896 4722
rect 2028 5754 1896 5822
rect 2028 5094 1896 5162
rect 2028 5534 1896 5602
rect 2028 5314 1896 5382
rect 2028 4874 1896 4942
rect 2028 4654 1896 4722
rect 2028 5754 1896 5822
rect 2028 5094 1896 5162
rect 2028 5534 1896 5602
rect 2028 5314 1896 5382
rect 2028 4874 1896 4942
rect 2028 10606 1896 10674
rect 2028 11706 1896 11774
rect 2028 11046 1896 11114
rect 2028 11486 1896 11554
rect 2028 11266 1896 11334
rect 2028 10826 1896 10894
rect 2028 10606 1896 10674
rect 2028 11706 1896 11774
rect 2028 11046 1896 11114
rect 2028 11486 1896 11554
rect 2028 11266 1896 11334
rect 2028 10826 1896 10894
rect 2028 10606 1896 10674
rect 2028 11706 1896 11774
rect 2028 11046 1896 11114
rect 2028 11486 1896 11554
rect 2028 11266 1896 11334
rect 2028 10826 1896 10894
rect 2028 10606 1896 10674
rect 2028 11706 1896 11774
rect 2028 11046 1896 11114
rect 2028 11486 1896 11554
rect 2028 11266 1896 11334
rect 2028 10826 1896 10894
rect 2028 10606 1896 10674
rect 2028 11706 1896 11774
rect 2028 11046 1896 11114
rect 2028 11486 1896 11554
rect 2028 11266 1896 11334
rect 2028 10826 1896 10894
rect 2028 10606 1896 10674
rect 2028 11706 1896 11774
rect 2028 11046 1896 11114
rect 2028 11486 1896 11554
rect 2028 11266 1896 11334
rect 2028 10826 1896 10894
rect 2028 190 1740 258
rect 2028 1290 1740 1358
rect 2028 630 1740 698
rect 2028 1070 1740 1138
rect 2028 850 1740 918
rect 2028 410 1740 478
rect 2028 190 1740 258
rect 2028 1290 1740 1358
rect 2028 630 1740 698
rect 2028 1070 1740 1138
rect 2028 850 1740 918
rect 2028 410 1740 478
rect 2028 190 1740 258
rect 2028 1290 1740 1358
rect 2028 630 1740 698
rect 2028 1070 1740 1138
rect 2028 850 1740 918
rect 2028 410 1740 478
rect 2028 190 1740 258
rect 2028 1290 1740 1358
rect 2028 630 1740 698
rect 2028 1070 1740 1138
rect 2028 850 1740 918
rect 2028 410 1740 478
rect 2028 190 1740 258
rect 2028 1290 1740 1358
rect 2028 630 1740 698
rect 2028 1070 1740 1138
rect 2028 850 1740 918
rect 2028 410 1740 478
rect 2028 190 1740 258
rect 2028 1290 1740 1358
rect 2028 630 1740 698
rect 2028 1070 1740 1138
rect 2028 850 1740 918
rect 2028 410 1740 478
rect 2028 6142 1740 6210
rect 2028 7242 1740 7310
rect 2028 6582 1740 6650
rect 2028 7022 1740 7090
rect 2028 6802 1740 6870
rect 2028 6362 1740 6430
rect 2028 6142 1740 6210
rect 2028 7242 1740 7310
rect 2028 6582 1740 6650
rect 2028 7022 1740 7090
rect 2028 6802 1740 6870
rect 2028 6362 1740 6430
rect 2028 6142 1740 6210
rect 2028 7242 1740 7310
rect 2028 6582 1740 6650
rect 2028 7022 1740 7090
rect 2028 6802 1740 6870
rect 2028 6362 1740 6430
rect 2028 6142 1740 6210
rect 2028 7242 1740 7310
rect 2028 6582 1740 6650
rect 2028 7022 1740 7090
rect 2028 6802 1740 6870
rect 2028 6362 1740 6430
rect 2028 6142 1740 6210
rect 2028 7242 1740 7310
rect 2028 6582 1740 6650
rect 2028 7022 1740 7090
rect 2028 6802 1740 6870
rect 2028 6362 1740 6430
rect 2028 6142 1740 6210
rect 2028 7242 1740 7310
rect 2028 6582 1740 6650
rect 2028 7022 1740 7090
rect 2028 6802 1740 6870
rect 2028 6362 1740 6430
rect 2028 9118 1584 9186
rect 2028 10218 1584 10286
rect 2028 9558 1584 9626
rect 2028 9998 1584 10066
rect 2028 9778 1584 9846
rect 2028 9338 1584 9406
rect 2028 9118 1584 9186
rect 2028 10218 1584 10286
rect 2028 9558 1584 9626
rect 2028 9998 1584 10066
rect 2028 9778 1584 9846
rect 2028 9338 1584 9406
rect 2028 9118 1584 9186
rect 2028 10218 1584 10286
rect 2028 9558 1584 9626
rect 2028 9998 1584 10066
rect 2028 9778 1584 9846
rect 2028 9338 1584 9406
rect 2028 9118 1584 9186
rect 2028 10218 1584 10286
rect 2028 9558 1584 9626
rect 2028 9998 1584 10066
rect 2028 9778 1584 9846
rect 2028 9338 1584 9406
rect 2028 9118 1584 9186
rect 2028 10218 1584 10286
rect 2028 9558 1584 9626
rect 2028 9998 1584 10066
rect 2028 9778 1584 9846
rect 2028 9338 1584 9406
rect 2028 9118 1584 9186
rect 2028 10218 1584 10286
rect 2028 9558 1584 9626
rect 2028 9998 1584 10066
rect 2028 9778 1584 9846
rect 2028 9338 1584 9406
rect 2028 1678 1428 1746
rect 2028 2778 1428 2846
rect 2028 2118 1428 2186
rect 2028 2558 1428 2626
rect 2028 2338 1428 2406
rect 2028 1898 1428 1966
rect 2028 1678 1428 1746
rect 2028 2778 1428 2846
rect 2028 2118 1428 2186
rect 2028 2558 1428 2626
rect 2028 2338 1428 2406
rect 2028 1898 1428 1966
rect 2028 1678 1428 1746
rect 2028 2778 1428 2846
rect 2028 2118 1428 2186
rect 2028 2558 1428 2626
rect 2028 2338 1428 2406
rect 2028 1898 1428 1966
rect 2028 1678 1428 1746
rect 2028 2778 1428 2846
rect 2028 2118 1428 2186
rect 2028 2558 1428 2626
rect 2028 2338 1428 2406
rect 2028 1898 1428 1966
rect 2028 1678 1428 1746
rect 2028 2778 1428 2846
rect 2028 2118 1428 2186
rect 2028 2558 1428 2626
rect 2028 2338 1428 2406
rect 2028 1898 1428 1966
rect 2028 1678 1428 1746
rect 2028 2778 1428 2846
rect 2028 2118 1428 2186
rect 2028 2558 1428 2626
rect 2028 2338 1428 2406
rect 2028 1898 1428 1966
rect 2028 3386 1272 3454
rect 2028 7850 1116 7918
rect 2028 7630 960 7698
rect 2028 8730 960 8798
rect 2028 8070 960 8138
rect 2028 8510 960 8578
rect 2028 7630 960 7698
rect 2028 8730 960 8798
rect 2028 8070 960 8138
rect 2028 8510 960 8578
rect 2028 7630 960 7698
rect 2028 8730 960 8798
rect 2028 8070 960 8138
rect 2028 8510 960 8578
rect 2028 7630 960 7698
rect 2028 8730 960 8798
rect 2028 8070 960 8138
rect 2028 8510 960 8578
rect 2028 8290 804 8358
rect 2028 3826 648 3894
rect 2028 4046 492 4114
rect 2028 3606 336 3674
rect 2028 4266 180 4334
use CAP32C_CV XC1
transform 1 0 2028 0 1 0
box 2028 0 10988 1488
use CAP32C_CV XC64a<0>
transform 1 0 2028 0 1 1488
box 2028 1488 10988 2976
use CAP32C_CV XC32a<0>
transform 1 0 2028 0 1 2976
box 2028 2976 10988 4464
use CAP32C_CV XC128a<1>
transform 1 0 2028 0 1 4464
box 2028 4464 10988 5952
use CAP32C_CV XC128b<2>
transform 1 0 2028 0 1 5952
box 2028 5952 10988 7440
use CAP32C_CV X16ab
transform 1 0 2028 0 1 7440
box 2028 7440 10988 8928
use CAP32C_CV XC64b<1>
transform 1 0 2028 0 1 8928
box 2028 8928 10988 10416
use CAP32C_CV XC0
transform 1 0 2028 0 1 10416
box 2028 10416 10988 11904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4654
box 2028 4654 2212 4722
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4596
box 1832 4596 1900 4780
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5754
box 2028 5754 2212 5822
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5696
box 1832 5696 1900 5880
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5094
box 2028 5094 2212 5162
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5036
box 1832 5036 1900 5220
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5534
box 2028 5534 2212 5602
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5476
box 1832 5476 1900 5660
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5314
box 2028 5314 2212 5382
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5256
box 1832 5256 1900 5440
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4874
box 2028 4874 2212 4942
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4816
box 1832 4816 1900 5000
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4654
box 2028 4654 2212 4722
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4596
box 1832 4596 1900 4780
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5754
box 2028 5754 2212 5822
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5696
box 1832 5696 1900 5880
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5094
box 2028 5094 2212 5162
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5036
box 1832 5036 1900 5220
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5534
box 2028 5534 2212 5602
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5476
box 1832 5476 1900 5660
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5314
box 2028 5314 2212 5382
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5256
box 1832 5256 1900 5440
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4874
box 2028 4874 2212 4942
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4816
box 1832 4816 1900 5000
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4654
box 2028 4654 2212 4722
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4596
box 1832 4596 1900 4780
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5754
box 2028 5754 2212 5822
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5696
box 1832 5696 1900 5880
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5094
box 2028 5094 2212 5162
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5036
box 1832 5036 1900 5220
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5534
box 2028 5534 2212 5602
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5476
box 1832 5476 1900 5660
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5314
box 2028 5314 2212 5382
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5256
box 1832 5256 1900 5440
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4874
box 2028 4874 2212 4942
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4816
box 1832 4816 1900 5000
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4654
box 2028 4654 2212 4722
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4596
box 1832 4596 1900 4780
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5754
box 2028 5754 2212 5822
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5696
box 1832 5696 1900 5880
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5094
box 2028 5094 2212 5162
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5036
box 1832 5036 1900 5220
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5534
box 2028 5534 2212 5602
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5476
box 1832 5476 1900 5660
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5314
box 2028 5314 2212 5382
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5256
box 1832 5256 1900 5440
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4874
box 2028 4874 2212 4942
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4816
box 1832 4816 1900 5000
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4654
box 2028 4654 2212 4722
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4596
box 1832 4596 1900 4780
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5754
box 2028 5754 2212 5822
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5696
box 1832 5696 1900 5880
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5094
box 2028 5094 2212 5162
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5036
box 1832 5036 1900 5220
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5534
box 2028 5534 2212 5602
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5476
box 1832 5476 1900 5660
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5314
box 2028 5314 2212 5382
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5256
box 1832 5256 1900 5440
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4874
box 2028 4874 2212 4942
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4816
box 1832 4816 1900 5000
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4654
box 2028 4654 2212 4722
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4596
box 1832 4596 1900 4780
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5754
box 2028 5754 2212 5822
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5696
box 1832 5696 1900 5880
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5094
box 2028 5094 2212 5162
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5036
box 1832 5036 1900 5220
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5534
box 2028 5534 2212 5602
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5476
box 1832 5476 1900 5660
use cut_M1M3_2x1 
transform 1 0 2028 0 1 5314
box 2028 5314 2212 5382
use cut_M2M3_1x2 
transform 1 0 1832 0 1 5256
box 1832 5256 1900 5440
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4874
box 2028 4874 2212 4942
use cut_M2M3_1x2 
transform 1 0 1832 0 1 4816
box 1832 4816 1900 5000
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10606
box 2028 10606 2212 10674
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10548
box 1832 10548 1900 10732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11706
box 2028 11706 2212 11774
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11648
box 1832 11648 1900 11832
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11046
box 2028 11046 2212 11114
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10988
box 1832 10988 1900 11172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11486
box 2028 11486 2212 11554
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11428
box 1832 11428 1900 11612
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11266
box 2028 11266 2212 11334
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11208
box 1832 11208 1900 11392
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10826
box 2028 10826 2212 10894
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10768
box 1832 10768 1900 10952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10606
box 2028 10606 2212 10674
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10548
box 1832 10548 1900 10732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11706
box 2028 11706 2212 11774
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11648
box 1832 11648 1900 11832
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11046
box 2028 11046 2212 11114
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10988
box 1832 10988 1900 11172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11486
box 2028 11486 2212 11554
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11428
box 1832 11428 1900 11612
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11266
box 2028 11266 2212 11334
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11208
box 1832 11208 1900 11392
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10826
box 2028 10826 2212 10894
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10768
box 1832 10768 1900 10952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10606
box 2028 10606 2212 10674
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10548
box 1832 10548 1900 10732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11706
box 2028 11706 2212 11774
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11648
box 1832 11648 1900 11832
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11046
box 2028 11046 2212 11114
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10988
box 1832 10988 1900 11172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11486
box 2028 11486 2212 11554
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11428
box 1832 11428 1900 11612
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11266
box 2028 11266 2212 11334
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11208
box 1832 11208 1900 11392
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10826
box 2028 10826 2212 10894
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10768
box 1832 10768 1900 10952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10606
box 2028 10606 2212 10674
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10548
box 1832 10548 1900 10732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11706
box 2028 11706 2212 11774
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11648
box 1832 11648 1900 11832
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11046
box 2028 11046 2212 11114
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10988
box 1832 10988 1900 11172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11486
box 2028 11486 2212 11554
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11428
box 1832 11428 1900 11612
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11266
box 2028 11266 2212 11334
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11208
box 1832 11208 1900 11392
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10826
box 2028 10826 2212 10894
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10768
box 1832 10768 1900 10952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10606
box 2028 10606 2212 10674
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10548
box 1832 10548 1900 10732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11706
box 2028 11706 2212 11774
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11648
box 1832 11648 1900 11832
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11046
box 2028 11046 2212 11114
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10988
box 1832 10988 1900 11172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11486
box 2028 11486 2212 11554
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11428
box 1832 11428 1900 11612
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11266
box 2028 11266 2212 11334
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11208
box 1832 11208 1900 11392
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10826
box 2028 10826 2212 10894
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10768
box 1832 10768 1900 10952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10606
box 2028 10606 2212 10674
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10548
box 1832 10548 1900 10732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11706
box 2028 11706 2212 11774
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11648
box 1832 11648 1900 11832
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11046
box 2028 11046 2212 11114
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10988
box 1832 10988 1900 11172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11486
box 2028 11486 2212 11554
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11428
box 1832 11428 1900 11612
use cut_M1M3_2x1 
transform 1 0 2028 0 1 11266
box 2028 11266 2212 11334
use cut_M2M3_1x2 
transform 1 0 1832 0 1 11208
box 1832 11208 1900 11392
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10826
box 2028 10826 2212 10894
use cut_M2M3_1x2 
transform 1 0 1832 0 1 10768
box 1832 10768 1900 10952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 190
box 2028 190 2212 258
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 316
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1290
box 2028 1290 2212 1358
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1232
box 1676 1232 1744 1416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 630
box 2028 630 2212 698
use cut_M2M3_1x2 
transform 1 0 1676 0 1 572
box 1676 572 1744 756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1070
box 2028 1070 2212 1138
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1012
box 1676 1012 1744 1196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 850
box 2028 850 2212 918
use cut_M2M3_1x2 
transform 1 0 1676 0 1 792
box 1676 792 1744 976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 410
box 2028 410 2212 478
use cut_M2M3_1x2 
transform 1 0 1676 0 1 352
box 1676 352 1744 536
use cut_M1M3_2x1 
transform 1 0 2028 0 1 190
box 2028 190 2212 258
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 316
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1290
box 2028 1290 2212 1358
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1232
box 1676 1232 1744 1416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 630
box 2028 630 2212 698
use cut_M2M3_1x2 
transform 1 0 1676 0 1 572
box 1676 572 1744 756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1070
box 2028 1070 2212 1138
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1012
box 1676 1012 1744 1196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 850
box 2028 850 2212 918
use cut_M2M3_1x2 
transform 1 0 1676 0 1 792
box 1676 792 1744 976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 410
box 2028 410 2212 478
use cut_M2M3_1x2 
transform 1 0 1676 0 1 352
box 1676 352 1744 536
use cut_M1M3_2x1 
transform 1 0 2028 0 1 190
box 2028 190 2212 258
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 316
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1290
box 2028 1290 2212 1358
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1232
box 1676 1232 1744 1416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 630
box 2028 630 2212 698
use cut_M2M3_1x2 
transform 1 0 1676 0 1 572
box 1676 572 1744 756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1070
box 2028 1070 2212 1138
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1012
box 1676 1012 1744 1196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 850
box 2028 850 2212 918
use cut_M2M3_1x2 
transform 1 0 1676 0 1 792
box 1676 792 1744 976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 410
box 2028 410 2212 478
use cut_M2M3_1x2 
transform 1 0 1676 0 1 352
box 1676 352 1744 536
use cut_M1M3_2x1 
transform 1 0 2028 0 1 190
box 2028 190 2212 258
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 316
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1290
box 2028 1290 2212 1358
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1232
box 1676 1232 1744 1416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 630
box 2028 630 2212 698
use cut_M2M3_1x2 
transform 1 0 1676 0 1 572
box 1676 572 1744 756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1070
box 2028 1070 2212 1138
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1012
box 1676 1012 1744 1196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 850
box 2028 850 2212 918
use cut_M2M3_1x2 
transform 1 0 1676 0 1 792
box 1676 792 1744 976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 410
box 2028 410 2212 478
use cut_M2M3_1x2 
transform 1 0 1676 0 1 352
box 1676 352 1744 536
use cut_M1M3_2x1 
transform 1 0 2028 0 1 190
box 2028 190 2212 258
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 316
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1290
box 2028 1290 2212 1358
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1232
box 1676 1232 1744 1416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 630
box 2028 630 2212 698
use cut_M2M3_1x2 
transform 1 0 1676 0 1 572
box 1676 572 1744 756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1070
box 2028 1070 2212 1138
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1012
box 1676 1012 1744 1196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 850
box 2028 850 2212 918
use cut_M2M3_1x2 
transform 1 0 1676 0 1 792
box 1676 792 1744 976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 410
box 2028 410 2212 478
use cut_M2M3_1x2 
transform 1 0 1676 0 1 352
box 1676 352 1744 536
use cut_M1M3_2x1 
transform 1 0 2028 0 1 190
box 2028 190 2212 258
use cut_M2M3_1x2 
transform 1 0 1676 0 1 132
box 1676 132 1744 316
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1290
box 2028 1290 2212 1358
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1232
box 1676 1232 1744 1416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 630
box 2028 630 2212 698
use cut_M2M3_1x2 
transform 1 0 1676 0 1 572
box 1676 572 1744 756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1070
box 2028 1070 2212 1138
use cut_M2M3_1x2 
transform 1 0 1676 0 1 1012
box 1676 1012 1744 1196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 850
box 2028 850 2212 918
use cut_M2M3_1x2 
transform 1 0 1676 0 1 792
box 1676 792 1744 976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 410
box 2028 410 2212 478
use cut_M2M3_1x2 
transform 1 0 1676 0 1 352
box 1676 352 1744 536
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6142
box 2028 6142 2212 6210
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6084
box 1676 6084 1744 6268
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7242
box 2028 7242 2212 7310
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7184
box 1676 7184 1744 7368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6582
box 2028 6582 2212 6650
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6524
box 1676 6524 1744 6708
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7022
box 2028 7022 2212 7090
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6964
box 1676 6964 1744 7148
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6802
box 2028 6802 2212 6870
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6744
box 1676 6744 1744 6928
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6362
box 2028 6362 2212 6430
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6304
box 1676 6304 1744 6488
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6142
box 2028 6142 2212 6210
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6084
box 1676 6084 1744 6268
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7242
box 2028 7242 2212 7310
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7184
box 1676 7184 1744 7368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6582
box 2028 6582 2212 6650
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6524
box 1676 6524 1744 6708
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7022
box 2028 7022 2212 7090
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6964
box 1676 6964 1744 7148
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6802
box 2028 6802 2212 6870
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6744
box 1676 6744 1744 6928
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6362
box 2028 6362 2212 6430
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6304
box 1676 6304 1744 6488
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6142
box 2028 6142 2212 6210
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6084
box 1676 6084 1744 6268
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7242
box 2028 7242 2212 7310
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7184
box 1676 7184 1744 7368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6582
box 2028 6582 2212 6650
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6524
box 1676 6524 1744 6708
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7022
box 2028 7022 2212 7090
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6964
box 1676 6964 1744 7148
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6802
box 2028 6802 2212 6870
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6744
box 1676 6744 1744 6928
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6362
box 2028 6362 2212 6430
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6304
box 1676 6304 1744 6488
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6142
box 2028 6142 2212 6210
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6084
box 1676 6084 1744 6268
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7242
box 2028 7242 2212 7310
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7184
box 1676 7184 1744 7368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6582
box 2028 6582 2212 6650
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6524
box 1676 6524 1744 6708
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7022
box 2028 7022 2212 7090
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6964
box 1676 6964 1744 7148
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6802
box 2028 6802 2212 6870
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6744
box 1676 6744 1744 6928
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6362
box 2028 6362 2212 6430
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6304
box 1676 6304 1744 6488
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6142
box 2028 6142 2212 6210
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6084
box 1676 6084 1744 6268
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7242
box 2028 7242 2212 7310
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7184
box 1676 7184 1744 7368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6582
box 2028 6582 2212 6650
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6524
box 1676 6524 1744 6708
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7022
box 2028 7022 2212 7090
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6964
box 1676 6964 1744 7148
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6802
box 2028 6802 2212 6870
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6744
box 1676 6744 1744 6928
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6362
box 2028 6362 2212 6430
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6304
box 1676 6304 1744 6488
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6142
box 2028 6142 2212 6210
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6084
box 1676 6084 1744 6268
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7242
box 2028 7242 2212 7310
use cut_M2M3_1x2 
transform 1 0 1676 0 1 7184
box 1676 7184 1744 7368
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6582
box 2028 6582 2212 6650
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6524
box 1676 6524 1744 6708
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7022
box 2028 7022 2212 7090
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6964
box 1676 6964 1744 7148
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6802
box 2028 6802 2212 6870
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6744
box 1676 6744 1744 6928
use cut_M1M3_2x1 
transform 1 0 2028 0 1 6362
box 2028 6362 2212 6430
use cut_M2M3_1x2 
transform 1 0 1676 0 1 6304
box 1676 6304 1744 6488
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9118
box 2028 9118 2212 9186
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9060
box 1520 9060 1588 9244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10218
box 2028 10218 2212 10286
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10160
box 1520 10160 1588 10344
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9558
box 2028 9558 2212 9626
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9500
box 1520 9500 1588 9684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9998
box 2028 9998 2212 10066
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9940
box 1520 9940 1588 10124
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9778
box 2028 9778 2212 9846
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9720
box 1520 9720 1588 9904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9338
box 2028 9338 2212 9406
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9280
box 1520 9280 1588 9464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9118
box 2028 9118 2212 9186
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9060
box 1520 9060 1588 9244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10218
box 2028 10218 2212 10286
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10160
box 1520 10160 1588 10344
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9558
box 2028 9558 2212 9626
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9500
box 1520 9500 1588 9684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9998
box 2028 9998 2212 10066
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9940
box 1520 9940 1588 10124
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9778
box 2028 9778 2212 9846
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9720
box 1520 9720 1588 9904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9338
box 2028 9338 2212 9406
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9280
box 1520 9280 1588 9464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9118
box 2028 9118 2212 9186
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9060
box 1520 9060 1588 9244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10218
box 2028 10218 2212 10286
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10160
box 1520 10160 1588 10344
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9558
box 2028 9558 2212 9626
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9500
box 1520 9500 1588 9684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9998
box 2028 9998 2212 10066
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9940
box 1520 9940 1588 10124
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9778
box 2028 9778 2212 9846
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9720
box 1520 9720 1588 9904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9338
box 2028 9338 2212 9406
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9280
box 1520 9280 1588 9464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9118
box 2028 9118 2212 9186
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9060
box 1520 9060 1588 9244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10218
box 2028 10218 2212 10286
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10160
box 1520 10160 1588 10344
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9558
box 2028 9558 2212 9626
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9500
box 1520 9500 1588 9684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9998
box 2028 9998 2212 10066
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9940
box 1520 9940 1588 10124
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9778
box 2028 9778 2212 9846
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9720
box 1520 9720 1588 9904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9338
box 2028 9338 2212 9406
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9280
box 1520 9280 1588 9464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9118
box 2028 9118 2212 9186
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9060
box 1520 9060 1588 9244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10218
box 2028 10218 2212 10286
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10160
box 1520 10160 1588 10344
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9558
box 2028 9558 2212 9626
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9500
box 1520 9500 1588 9684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9998
box 2028 9998 2212 10066
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9940
box 1520 9940 1588 10124
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9778
box 2028 9778 2212 9846
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9720
box 1520 9720 1588 9904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9338
box 2028 9338 2212 9406
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9280
box 1520 9280 1588 9464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9118
box 2028 9118 2212 9186
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9060
box 1520 9060 1588 9244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 10218
box 2028 10218 2212 10286
use cut_M2M3_1x2 
transform 1 0 1520 0 1 10160
box 1520 10160 1588 10344
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9558
box 2028 9558 2212 9626
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9500
box 1520 9500 1588 9684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9998
box 2028 9998 2212 10066
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9940
box 1520 9940 1588 10124
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9778
box 2028 9778 2212 9846
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9720
box 1520 9720 1588 9904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 9338
box 2028 9338 2212 9406
use cut_M2M3_1x2 
transform 1 0 1520 0 1 9280
box 1520 9280 1588 9464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1678
box 2028 1678 2212 1746
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1620
box 1364 1620 1432 1804
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2778
box 2028 2778 2212 2846
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2720
box 1364 2720 1432 2904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2118
box 2028 2118 2212 2186
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2060
box 1364 2060 1432 2244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2558
box 2028 2558 2212 2626
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2500
box 1364 2500 1432 2684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2338
box 2028 2338 2212 2406
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2280
box 1364 2280 1432 2464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1898
box 2028 1898 2212 1966
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1840
box 1364 1840 1432 2024
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1678
box 2028 1678 2212 1746
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1620
box 1364 1620 1432 1804
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2778
box 2028 2778 2212 2846
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2720
box 1364 2720 1432 2904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2118
box 2028 2118 2212 2186
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2060
box 1364 2060 1432 2244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2558
box 2028 2558 2212 2626
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2500
box 1364 2500 1432 2684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2338
box 2028 2338 2212 2406
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2280
box 1364 2280 1432 2464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1898
box 2028 1898 2212 1966
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1840
box 1364 1840 1432 2024
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1678
box 2028 1678 2212 1746
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1620
box 1364 1620 1432 1804
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2778
box 2028 2778 2212 2846
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2720
box 1364 2720 1432 2904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2118
box 2028 2118 2212 2186
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2060
box 1364 2060 1432 2244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2558
box 2028 2558 2212 2626
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2500
box 1364 2500 1432 2684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2338
box 2028 2338 2212 2406
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2280
box 1364 2280 1432 2464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1898
box 2028 1898 2212 1966
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1840
box 1364 1840 1432 2024
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1678
box 2028 1678 2212 1746
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1620
box 1364 1620 1432 1804
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2778
box 2028 2778 2212 2846
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2720
box 1364 2720 1432 2904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2118
box 2028 2118 2212 2186
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2060
box 1364 2060 1432 2244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2558
box 2028 2558 2212 2626
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2500
box 1364 2500 1432 2684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2338
box 2028 2338 2212 2406
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2280
box 1364 2280 1432 2464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1898
box 2028 1898 2212 1966
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1840
box 1364 1840 1432 2024
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1678
box 2028 1678 2212 1746
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1620
box 1364 1620 1432 1804
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2778
box 2028 2778 2212 2846
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2720
box 1364 2720 1432 2904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2118
box 2028 2118 2212 2186
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2060
box 1364 2060 1432 2244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2558
box 2028 2558 2212 2626
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2500
box 1364 2500 1432 2684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2338
box 2028 2338 2212 2406
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2280
box 1364 2280 1432 2464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1898
box 2028 1898 2212 1966
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1840
box 1364 1840 1432 2024
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1678
box 2028 1678 2212 1746
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1620
box 1364 1620 1432 1804
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2778
box 2028 2778 2212 2846
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2720
box 1364 2720 1432 2904
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2118
box 2028 2118 2212 2186
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2060
box 1364 2060 1432 2244
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2558
box 2028 2558 2212 2626
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2500
box 1364 2500 1432 2684
use cut_M1M3_2x1 
transform 1 0 2028 0 1 2338
box 2028 2338 2212 2406
use cut_M2M3_1x2 
transform 1 0 1364 0 1 2280
box 1364 2280 1432 2464
use cut_M1M3_2x1 
transform 1 0 2028 0 1 1898
box 2028 1898 2212 1966
use cut_M2M3_1x2 
transform 1 0 1364 0 1 1840
box 1364 1840 1432 2024
use cut_M1M3_2x1 
transform 1 0 2028 0 1 3386
box 2028 3386 2212 3454
use cut_M2M3_1x2 
transform 1 0 1208 0 1 3328
box 1208 3328 1276 3512
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7850
box 2028 7850 2212 7918
use cut_M2M3_1x2 
transform 1 0 1052 0 1 7792
box 1052 7792 1120 7976
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7630
box 2028 7630 2212 7698
use cut_M2M3_1x2 
transform 1 0 896 0 1 7572
box 896 7572 964 7756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8730
box 2028 8730 2212 8798
use cut_M2M3_1x2 
transform 1 0 896 0 1 8672
box 896 8672 964 8856
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8070
box 2028 8070 2212 8138
use cut_M2M3_1x2 
transform 1 0 896 0 1 8012
box 896 8012 964 8196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8510
box 2028 8510 2212 8578
use cut_M2M3_1x2 
transform 1 0 896 0 1 8452
box 896 8452 964 8636
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7630
box 2028 7630 2212 7698
use cut_M2M3_1x2 
transform 1 0 896 0 1 7572
box 896 7572 964 7756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8730
box 2028 8730 2212 8798
use cut_M2M3_1x2 
transform 1 0 896 0 1 8672
box 896 8672 964 8856
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8070
box 2028 8070 2212 8138
use cut_M2M3_1x2 
transform 1 0 896 0 1 8012
box 896 8012 964 8196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8510
box 2028 8510 2212 8578
use cut_M2M3_1x2 
transform 1 0 896 0 1 8452
box 896 8452 964 8636
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7630
box 2028 7630 2212 7698
use cut_M2M3_1x2 
transform 1 0 896 0 1 7572
box 896 7572 964 7756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8730
box 2028 8730 2212 8798
use cut_M2M3_1x2 
transform 1 0 896 0 1 8672
box 896 8672 964 8856
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8070
box 2028 8070 2212 8138
use cut_M2M3_1x2 
transform 1 0 896 0 1 8012
box 896 8012 964 8196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8510
box 2028 8510 2212 8578
use cut_M2M3_1x2 
transform 1 0 896 0 1 8452
box 896 8452 964 8636
use cut_M1M3_2x1 
transform 1 0 2028 0 1 7630
box 2028 7630 2212 7698
use cut_M2M3_1x2 
transform 1 0 896 0 1 7572
box 896 7572 964 7756
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8730
box 2028 8730 2212 8798
use cut_M2M3_1x2 
transform 1 0 896 0 1 8672
box 896 8672 964 8856
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8070
box 2028 8070 2212 8138
use cut_M2M3_1x2 
transform 1 0 896 0 1 8012
box 896 8012 964 8196
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8510
box 2028 8510 2212 8578
use cut_M2M3_1x2 
transform 1 0 896 0 1 8452
box 896 8452 964 8636
use cut_M1M3_2x1 
transform 1 0 2028 0 1 8290
box 2028 8290 2212 8358
use cut_M2M3_1x2 
transform 1 0 740 0 1 8232
box 740 8232 808 8416
use cut_M1M3_2x1 
transform 1 0 2028 0 1 3826
box 2028 3826 2212 3894
use cut_M2M3_1x2 
transform 1 0 584 0 1 3768
box 584 3768 652 3952
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4046
box 2028 4046 2212 4114
use cut_M2M3_1x2 
transform 1 0 428 0 1 3988
box 428 3988 496 4172
use cut_M1M3_2x1 
transform 1 0 2028 0 1 3606
box 2028 3606 2212 3674
use cut_M2M3_1x2 
transform 1 0 272 0 1 3548
box 272 3548 340 3732
use cut_M1M3_2x1 
transform 1 0 2028 0 1 4266
box 2028 4266 2212 4334
use cut_M2M3_1x2 
transform 1 0 116 0 1 4208
box 116 4208 184 4392
use cut_M1M2_1x2 
transform 1 0 2340 0 1 3108
box 2340 3108 2408 3292
use cut_M1M2_1x2 
transform 1 0 2340 0 1 3108
box 2340 3108 2408 3292
<< labels >>
flabel m1 s 1836 4596 1896 11904 0 FreeSans 400 0 0 0 CP<11>
port 1 nsew
flabel m1 s 1680 132 1740 11904 0 FreeSans 400 0 0 0 CP<10>
port 2 nsew
flabel m1 s 1524 9060 1584 11904 0 FreeSans 400 0 0 0 CP<9>
port 3 nsew
flabel m1 s 1368 1620 1428 11904 0 FreeSans 400 0 0 0 CP<8>
port 4 nsew
flabel m1 s 1212 3328 1272 11904 0 FreeSans 400 0 0 0 CP<7>
port 5 nsew
flabel m1 s 1056 7792 1116 11904 0 FreeSans 400 0 0 0 CP<6>
port 6 nsew
flabel m1 s 900 7572 960 11904 0 FreeSans 400 0 0 0 CP<5>
port 7 nsew
flabel m1 s 744 8232 804 11904 0 FreeSans 400 0 0 0 CP<4>
port 8 nsew
flabel m1 s 588 3768 648 11904 0 FreeSans 400 0 0 0 CP<3>
port 9 nsew
flabel m1 s 432 3988 492 11904 0 FreeSans 400 0 0 0 CP<2>
port 10 nsew
flabel m1 s 276 3548 336 11904 0 FreeSans 400 0 0 0 CP<1>
port 11 nsew
flabel m1 s 120 4208 180 11904 0 FreeSans 400 0 0 0 CP<0>
port 12 nsew
flabel m1 s 2340 0 10920 68 0 FreeSans 400 0 0 0 AVSS
port 13 nsew
flabel m3 s 2340 10416 2408 11964 0 FreeSans 400 0 0 0 CTOP
port 14 nsew
<< end >>
