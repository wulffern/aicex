magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 1280
<< locali >>
rect 720 1170 874 1230
rect 874 50 1380 110
rect 874 1170 1380 1230
rect 874 50 934 1230
rect 330 130 390 1150
rect 1710 130 1770 510
rect 1710 770 1770 1150
rect 690 210 750 430
rect 690 530 750 750
rect 690 850 750 1070
rect 1350 210 1410 430
rect 1350 530 1410 750
rect 1350 850 1410 1070
rect 1650 130 1830 190
rect 1650 770 1830 830
rect 270 450 450 510
rect 630 1170 810 1230
<< m3 >>
rect 1290 0 1474 1280
rect 630 0 814 1280
rect 1290 0 1474 1280
rect 630 0 814 1280
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1050 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1050 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1050 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1050 1280
use PCHDL MP0
transform 1 0 1050 0 1 0
box 1050 0 2100 320
use PCHDL MP1
transform 1 0 1050 0 1 320
box 1050 320 2100 640
use PCHDL MP2
transform 1 0 1050 0 1 640
box 1050 640 2100 960
use PCHDL MP3
transform 1 0 1050 0 1 960
box 1050 960 2100 1280
use cut_M1M4_2x1 
transform 1 0 1290 0 1 530
box 1290 530 1474 598
use cut_M1M4_2x1 
transform 1 0 1290 0 1 690
box 1290 690 1474 758
use cut_M1M4_2x1 
transform 1 0 630 0 1 50
box 630 50 814 118
use cut_M1M4_2x1 
transform 1 0 630 0 1 530
box 630 530 814 598
use cut_M1M4_2x1 
transform 1 0 630 0 1 690
box 630 690 814 758
<< labels >>
flabel locali s 1650 130 1830 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 1650 770 1830 830 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 270 450 450 510 0 FreeSans 400 0 0 0 RST
port 3 nsew
flabel locali s 630 1170 810 1230 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel m3 s 1290 0 1474 1280 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 630 0 814 1280 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
