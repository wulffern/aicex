magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 640
<< locali >>
rect 800 210 968 270
rect 800 370 968 430
rect 968 210 1520 270
rect 968 370 1520 430
rect 968 210 1028 430
rect 370 130 430 510
rect 1890 130 1950 510
<< poly >>
rect 280 142 2040 178
rect 280 462 2040 498
<< m3 >>
rect 1400 0 1600 640
rect 680 0 880 640
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use cut_M1M4_2x1 
transform 1 0 1400 0 1 50
box 1400 50 1600 118
use cut_M1M4_2x1 
transform 1 0 1400 0 1 530
box 1400 530 1600 598
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
use cut_M1M4_2x1 
transform 1 0 680 0 1 530
box 680 530 880 598
<< labels >>
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 A
port 1 nsew
flabel locali s 680 210 920 270 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel locali s 2200 120 2440 200 0 FreeSans 400 0 0 0 BULKP
port 3 nsew
flabel locali s -120 120 120 200 0 FreeSans 400 0 0 0 BULKN
port 4 nsew
flabel m3 s 1400 0 1600 640 0 FreeSans 400 0 0 0 AVDD
port 5 nsew
flabel m3 s 680 0 880 640 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
<< end >>
