
*-------------------------------------------------------------
* SUNTR_PCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDL D G S B
XMM1 D G S B sky130_fd_pr__pfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDL <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDL D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLR D G S B
XMM1 D G S B sky130_fd_pr__nfet_01v8  l=0.18  nf=1  w=1.08  
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLCM D G S B
XM0 N0 G S B SUNTR_NCHDL
XM1 N1 G N0 B SUNTR_NCHDL
XM2 N2 G N1 B SUNTR_NCHDL
XM3 N3 G N2 B SUNTR_NCHDL
XM4 N4 G N3 B SUNTR_NCHDL
XM5 N5 G N4 B SUNTR_NCHDL
XM6 N6 G N5 B SUNTR_NCHDL
XM7 N7 G N6 B SUNTR_NCHDL
XM8 D G N7 B SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLCM <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLCM D G S B
XM0 N0 G S B SUNTR_PCHDL
XM7 D G N0 B SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLA D G S B
XM0 D G S B SUNTR_NCHDL
XM1 S G D B SUNTR_NCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLA <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLA D G S B
XM0 D G S B SUNTR_PCHDL
XM1 S G D B SUNTR_PCHDL
XM2 D G S B SUNTR_PCHDL
XM3 S G D B SUNTR_PCHDL
XM4 D G S B SUNTR_PCHDL
XM5 S G D B SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NCHDLCM2 D G S B
XM0 D G S B SUNTR_NCHDLCM
XM1 S G D B SUNTR_NCHDLCM
.ENDS

*-------------------------------------------------------------
* SUNTR_PCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_PCHDLCM2 D G S B
XM0 D G S B SUNTR_PCHDLCM
XM1 S G D B SUNTR_PCHDLCM
.ENDS

*-------------------------------------------------------------
* SUNTR_CPCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_CPCHDLCM2 D G CG S CS B
XM0 CS G S B SUNTR_PCHDLCM2
XM1 D CG CS B SUNTR_PCHDLA
.ENDS

*-------------------------------------------------------------
* SUNTR_CNCHDLCM2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_CNCHDLCM2 D G CG S CS B
XM0 CS G S B SUNTR_NCHDLCM2
XM1 D CG CS B SUNTR_NCHDLA
.ENDS

*-------------------------------------------------------------
* SUNTR_RES12 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RES12 N P B
XRR1_0 N INT_0 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_1 INT_0 P B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
.ENDS

*-------------------------------------------------------------
* SUNTR_RES25 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RES25 N P B
XRR1_0 N INT_0 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_1 INT_0 INT_1 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_2 INT_1 INT_2 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_3 INT_2 P B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
.ENDS

*-------------------------------------------------------------
* SUNTR_RES100 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RES100 N P B
XRR1_0 N INT_0 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_1 INT_0 INT_1 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_2 INT_1 INT_2 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_3 INT_2 INT_3 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_4 INT_3 INT_4 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_5 INT_4 INT_5 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_6 INT_5 INT_6 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_7 INT_6 INT_7 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_8 INT_7 INT_8 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_9 INT_8 P B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
.ENDS

*-------------------------------------------------------------
* SUNTR_RES200 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RES200 N P B
XRR1_0 N INT_0 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_1 INT_0 INT_1 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_2 INT_1 INT_2 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_3 INT_2 INT_3 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_4 INT_3 INT_4 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_5 INT_4 INT_5 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_6 INT_5 INT_6 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_7 INT_6 INT_7 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_8 INT_7 INT_8 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_9 INT_8 INT_9 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_10 INT_9 INT_10 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_11 INT_10 INT_11 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_12 INT_11 INT_12 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_13 INT_12 INT_13 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_14 INT_13 INT_14 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_15 INT_14 INT_15 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_16 INT_15 INT_16 B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
XRR1_17 INT_16 P B sky130_fd_pr__res_high_po  l=8.8  w=0.54  
.ENDS

*-------------------------------------------------------------
* SUNTR_RPPO_12k <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RPPO_12k P N B
XA1 N P B SUNTR_RES12
.ENDS

*-------------------------------------------------------------
* SUNTR_RPPO_25k <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RPPO_25k P N B
XA1 N P B SUNTR_RES25
.ENDS

*-------------------------------------------------------------
* SUNTR_RPPO_100k <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RPPO_100k P N B
XA1 N P B SUNTR_RES100
.ENDS

*-------------------------------------------------------------
* SUNTR_RPPO_200k <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RPPO_200k P N B
XA1 N P B SUNTR_RES200
.ENDS

*-------------------------------------------------------------
* SUNTR_TAPCELLB_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TAPCELLB_CV AVDD AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTR_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_TIEH_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TIEH_CV Y AVDD AVSS
XMN0 A A AVSS AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_TIEL_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TIEL_CV Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMP0 A A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX1_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX2_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX4_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
XMP2 Y A AVDD AVDD SUNTR_PCHDL
XMP3 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVX8_CV A Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMN4 Y A AVSS AVSS SUNTR_NCHDL
XMN5 AVSS A Y AVSS SUNTR_NCHDL
XMN6 Y A AVSS AVSS SUNTR_NCHDL
XMN7 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD A Y AVDD SUNTR_PCHDL
XMP2 Y A AVDD AVDD SUNTR_PCHDL
XMP3 AVDD A Y AVDD SUNTR_PCHDL
XMP4 Y A AVDD AVDD SUNTR_PCHDL
XMP5 AVDD A Y AVDD SUNTR_PCHDL
XMP6 Y A AVDD AVDD SUNTR_PCHDL
XMP7 AVDD A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_BFX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_BFX1_CV A Y AVDD AVSS
XMN0 AVSS A B AVSS SUNTR_NCHDL
XMN1 Y B AVSS AVSS SUNTR_NCHDL
XMP0 AVDD A B AVDD SUNTR_PCHDL
XMP1 Y B AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NRX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NRX1_CV A B Y AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS B Y AVSS SUNTR_NCHDL
XMP0 N1 A AVDD AVDD SUNTR_PCHDL
XMP1 Y B N1 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NDX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NDX1_CV A B Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y B N1 AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD B Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_ORX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ORX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NRX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ORX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ORX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NRX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ORX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ORX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NRX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX1_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX2_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX4_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_ANX8_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_ANX8_CV A B Y AVDD AVSS
XA1 A B YN AVDD AVSS SUNTR_NDX1_CV
XA2 YN Y AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_DFTSPCX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFTSPCX1_CV D CK Q AVDD AVSS
XMN0 N1 D AVSS AVSS SUNTR_NCHDL
XMN2 N2 CK Q AVSS SUNTR_NCHDL
XMN1 AVSS N1 N2 AVSS SUNTR_NCHDL
XMP1 N3 D AVDD AVDD SUNTR_PCHDL
XMP0 N1 CK N3 AVDD SUNTR_PCHDL
XMP2 Q N1 AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_IVTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_IVTRIX1_CV A C CN Y AVDD AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y C N1 AVSS SUNTR_NCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NDTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NDTRIX1_CV A C CN RN Y AVDD AVSS
XMN2 N1 RN AVSS AVSS SUNTR_NCHDL
XMN0 N2 A N1 AVSS SUNTR_NCHDL
XMN1 Y C N2 AVSS SUNTR_NCHDL
XMP2 AVDD RN N2 AVDD SUNTR_PCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_NRTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_NRTRIX1_CV A C CN B Y AVDD AVSS
XMN2 N1 B AVSS AVSS SUNTR_NCHDL
XMN0 AVSS A N1 AVSS SUNTR_NCHDL
XMN1 N1 C Y AVSS SUNTR_NCHDL
XMP2 N2 B AVDD AVDD SUNTR_PCHDL
XMP0 AVDD A N2 AVDD SUNTR_PCHDL
XMP1 N2 CN Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_DFRNQNX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
XA0 AVDD AVSS SUNTR_TAPCELLB_CV
XA1 CK RN CKN AVDD AVSS SUNTR_NDX1_CV
XA2 CKN CKB AVDD AVSS SUNTR_IVX1_CV
XA3 D CKN CKB A0 AVDD AVSS SUNTR_IVTRIX1_CV
XA4 A1 CKB CKN A0 AVDD AVSS SUNTR_IVTRIX1_CV
XA5 A0 A1 AVDD AVSS SUNTR_IVX1_CV
XA6 A1 CKB CKN QN AVDD AVSS SUNTR_IVTRIX1_CV
XA7 Q CKN CKB RN QN AVDD AVSS SUNTR_NDTRIX1_CV
XA8 QN Q AVDD AVSS SUNTR_IVX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_SCX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SCX1_CV A Y AVDD AVSS
XA2 N1 A AVSS AVSS SUNTR_NCHDL
XA3 SCO A N1 AVSS SUNTR_NCHDL
XA4a AVDD SCO N1 AVSS SUNTR_NCHDL
XA4b AVDD SCO N1 AVSS SUNTR_NCHDL
XA5 Y SCO AVSS AVSS SUNTR_NCHDL
XB0 N2 A AVDD AVDD SUNTR_PCHDL
XB1 SCO A N2 AVDD SUNTR_PCHDL
XB3a N2 SCO AVSS AVDD SUNTR_PCHDL
XB3b N2 SCO AVSS AVDD SUNTR_PCHDL
XB4 Y SCO AVDD AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_SWX2_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SWX2_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A VREF AVDD SUNTR_PCHDL
XMP1 VREF A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_SWX4_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SWX4_CV A Y VREF AVDD AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS A Y AVSS SUNTR_NCHDL
XMN2 Y A AVSS AVSS SUNTR_NCHDL
XMN3 AVSS A Y AVSS SUNTR_NCHDL
XMP0 Y A VREF AVDD SUNTR_PCHDL
XMP1 VREF A Y AVDD SUNTR_PCHDL
XMP2 Y A VREF AVDD SUNTR_PCHDL
XMP3 VREF A Y AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_TGPD_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_TGPD_CV C A B AVDD AVSS
XMN0 AVSS C CN AVSS SUNTR_NCHDL
XMN1 B C AVSS AVSS SUNTR_NCHDL
XMN2 A CN B AVSS SUNTR_NCHDL
XMP0 AVDD C CN AVDD SUNTR_PCHDL
XMP1_DMY B AVDD AVDD AVDD SUNTR_PCHDL
XMP2 A C B AVDD SUNTR_PCHDL
.ENDS

*-------------------------------------------------------------
* SUNTR_DFTRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_DFTRIX1_CV D CK C CN Y AVDD AVSS
XA3 AVDD AVSS SUNTR_TAPCELLB_CV
XA2 D CK C NC QN AVDD AVSS SUNTR_DFRNQNX1_CV
XA0 QN C CN Y AVDD AVSS SUNTR_IVTRIX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_RG12TRIX1_CV <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_RG12TRIX1_CV D_11 D_10 D_9 D_8 D_7 D_6 D_5 D_4 D_3 D_2 D_1 D_0 CK C CN Y_11 Y_10 Y_9 Y_8 Y_7 Y_6 Y_5 Y_4 Y_3 Y_2 Y_1 Y_0 AVDD AVSS
XA0 D_11 CK C CN Y_11 AVDD AVSS SUNTR_DFTRIX1_CV
XB1 D_10 CK C CN Y_10 AVDD AVSS SUNTR_DFTRIX1_CV
XC2 D_9 CK C CN Y_9 AVDD AVSS SUNTR_DFTRIX1_CV
XD3 D_8 CK C CN Y_8 AVDD AVSS SUNTR_DFTRIX1_CV
XE4 D_7 CK C CN Y_7 AVDD AVSS SUNTR_DFTRIX1_CV
XF5 D_6 CK C CN Y_6 AVDD AVSS SUNTR_DFTRIX1_CV
XG6 D_5 CK C CN Y_5 AVDD AVSS SUNTR_DFTRIX1_CV
XH7 D_4 CK C CN Y_4 AVDD AVSS SUNTR_DFTRIX1_CV
XI8 D_3 CK C CN Y_3 AVDD AVSS SUNTR_DFTRIX1_CV
XJ9 D_2 CK C CN Y_2 AVDD AVSS SUNTR_DFTRIX1_CV
XK10 D_1 CK C CN Y_1 AVDD AVSS SUNTR_DFTRIX1_CV
XL11 D_0 CK C CN Y_0 AVDD AVSS SUNTR_DFTRIX1_CV
.ENDS

*-------------------------------------------------------------
* SUNTR_SUN_TR <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT SUNTR_SUN_TR AVDD AVSS
XA0 AVDD AVSS SUNTR_TAPCELLB_CV
XA1 Y1 AVDD AVSS SUNTR_TIEH_CV
XA2 Y2 AVDD AVSS SUNTR_TIEL_CV
XB0 AVDD AVSS SUNTR_TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS SUNTR_IVX1_CV
XB4 A4 Y4 AVDD AVSS SUNTR_IVX2_CV
XB5 A5 Y5 AVDD AVSS SUNTR_IVX4_CV
XB6 A6 Y6 AVDD AVSS SUNTR_IVX8_CV
XC0 AVDD AVSS SUNTR_TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS SUNTR_BFX1_CV
XD0 AVDD AVSS SUNTR_TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS SUNTR_NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS SUNTR_NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS SUNTR_ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS SUNTR_ANX1_CV
XE0 AVDD AVSS SUNTR_TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SUNTR_SCX1_CV
XF0 AVDD AVSS SUNTR_TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SUNTR_SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SUNTR_SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS SUNTR_TGPD_CV
.ENDS
