magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect 0 0 2100 10560
<< locali >>
rect 360 4610 514 4670
rect 514 4050 720 4110
rect 514 4050 574 4670
rect 360 5890 514 5950
rect 514 5330 720 5390
rect 514 5330 574 5950
rect 1526 3970 1740 4030
rect 1380 3730 1526 3790
rect 1526 3730 1586 4030
rect 360 8130 514 8190
rect 514 7890 720 7950
rect 514 7890 574 8190
rect 330 8130 390 8510
rect 390 9030 514 9090
rect 514 8850 720 8910
rect 514 8850 574 9090
rect 390 9090 450 9150
rect 390 9350 514 9410
rect 514 9170 720 9230
rect 514 9170 574 9410
rect 390 9410 450 9470
rect 360 10050 514 10110
rect 514 9650 720 9710
rect 514 9650 574 10110
rect 1380 5970 1534 6030
rect 1534 6530 1740 6590
rect 1534 5970 1594 6590
rect 1650 3650 1830 3710
rect 270 3010 450 3070
rect 270 9730 450 9790
rect 1290 10130 1470 10190
rect 270 6850 450 6910
rect 630 8210 810 8270
<< m1 >>
rect 360 5250 514 5310
rect 514 2770 720 2830
rect 514 2770 574 5318
rect 1740 7810 1894 7870
rect 1380 690 1894 750
rect 1894 690 1954 7878
rect 360 8770 514 8830
rect 514 7570 720 7630
rect 514 7570 574 8838
rect 1380 4690 1534 4750
rect 1534 7170 1740 7230
rect 1534 4690 1594 7238
<< m3 >>
rect 1828 4370 1896 6474
rect 266 4606 450 4674
rect 878 4628 946 4812
rect 1014 5268 1082 5452
rect 1150 5908 1218 6092
rect 1770 4370 1954 4554
rect 1290 0 1474 10560
rect 630 0 814 10560
rect 1290 0 1474 10560
rect 630 0 814 10560
<< m2 >>
rect 266 2046 450 2114
rect 266 446 450 514
rect 1286 686 1470 754
use DMY_CV XA0a
transform 1 0 0 0 1 0
box 0 0 0 0
use SARMRYX1_CV XA1
transform 1 0 0 0 1 0
box 0 0 2100 3840
use SWX2_CV XA2
transform 1 0 0 0 1 3840
box 0 3840 2100 4480
use SWX2_CV XA3
transform 1 0 0 0 1 4480
box 0 4480 2100 5120
use SWX2_CV XA4
transform 1 0 0 0 1 5120
box 0 5120 2100 5760
use SWX2_CV XA5
transform 1 0 0 0 1 5760
box 0 5760 2100 6400
use SARCEX1_CV XA6
transform 1 0 0 0 1 6400
box 0 6400 2100 7680
use IVX1_CV XA7
transform 1 0 0 0 1 7680
box 0 7680 2100 8000
use IVX1_CV XA8
transform 1 0 0 0 1 8000
box 0 8000 2100 8320
use NDX1_CV XA9
transform 1 0 0 0 1 8320
box 0 8320 2100 8960
use IVX1_CV XA10
transform 1 0 0 0 1 8960
box 0 8960 2100 9280
use NRX1_CV XA11
transform 1 0 0 0 1 9280
box 0 9280 2100 9920
use IVX1_CV XA12
transform 1 0 0 0 1 9920
box 0 9920 2100 10240
use TAPCELLB_CV XA13
transform 1 0 0 0 1 10240
box 0 10240 2100 10560
use DMY_CV XA14
transform 1 0 0 0 1 10560
box 0 10560 0 10560
use cut_M1M2_2x1 
transform 1 0 270 0 1 5250
box 270 5250 454 5318
use cut_M1M2_2x1 
transform 1 0 630 0 1 2770
box 630 2770 814 2838
use cut_M1M2_2x1 
transform 1 0 1650 0 1 7810
box 1650 7810 1834 7878
use cut_M1M2_2x1 
transform 1 0 1290 0 1 690
box 1290 690 1474 758
use cut_M1M2_2x1 
transform 1 0 270 0 1 8770
box 270 8770 454 8838
use cut_M1M2_2x1 
transform 1 0 630 0 1 7570
box 630 7570 814 7638
use cut_M1M2_2x1 
transform 1 0 1290 0 1 4690
box 1290 4690 1474 4758
use cut_M1M2_2x1 
transform 1 0 1650 0 1 7170
box 1650 7170 1834 7238
use cut_M1M4_2x1 
transform 1 0 266 0 1 4606
box 266 4606 450 4674
use cut_M1M4_1x2 
transform 1 0 878 0 1 4628
box 878 4628 946 4812
use cut_M1M4_1x2 
transform 1 0 1014 0 1 5268
box 1014 5268 1082 5452
use cut_M1M4_1x2 
transform 1 0 1150 0 1 5908
box 1150 5908 1218 6092
use cut_M2M3_2x1 
transform 1 0 1286 0 1 686
box 1286 686 1470 754
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 446
box 266 446 450 514
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
use cut_M2M3_2x1 
transform 1 0 266 0 1 2046
box 266 2046 450 2114
<< labels >>
flabel m2 s 266 2046 450 2114 0 FreeSans 400 0 0 0 CMP_OP
port 1 nsew
flabel locali s 1650 3650 1830 3710 0 FreeSans 400 0 0 0 RST_N
port 2 nsew
flabel m2 s 266 446 450 514 0 FreeSans 400 0 0 0 EN
port 3 nsew
flabel locali s 270 3010 450 3070 0 FreeSans 400 0 0 0 CMP_ON
port 4 nsew
flabel m2 s 1286 686 1470 754 0 FreeSans 400 0 0 0 ENO
port 5 nsew
flabel m3 s 266 4606 450 4674 0 FreeSans 400 0 0 0 CN1
port 6 nsew
flabel m3 s 878 4628 946 4812 0 FreeSans 400 0 0 0 CP1
port 7 nsew
flabel m3 s 1014 5268 1082 5452 0 FreeSans 400 0 0 0 CP0
port 8 nsew
flabel m3 s 1150 5908 1218 6092 0 FreeSans 400 0 0 0 CN0
port 9 nsew
flabel locali s 270 9730 450 9790 0 FreeSans 400 0 0 0 CEIN
port 10 nsew
flabel locali s 1290 10130 1470 10190 0 FreeSans 400 0 0 0 CEO
port 11 nsew
flabel locali s 270 6850 450 6910 0 FreeSans 400 0 0 0 CKS
port 12 nsew
flabel locali s 630 8210 810 8270 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 1770 4370 1954 4554 0 FreeSans 400 0 0 0 VREF
port 14 nsew
flabel m3 s 1290 0 1474 10560 0 FreeSans 400 0 0 0 AVDD
port 15 nsew
flabel m3 s 630 0 814 10560 0 FreeSans 400 0 0 0 AVSS
port 16 nsew
<< end >>
