magic
tech sky130A
magscale 1 2
timestamp 1659354040
<< checkpaint >>
rect 0 0 0 0
<< labels >>
<< end >>
