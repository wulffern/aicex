magic
tech sky130A
magscale 1 2
timestamp 1664575200
<< checkpaint >>
rect 0 0 1260 528
<< pdiff >>
rect 288 132 504 220
rect 288 220 504 308
rect 288 308 504 396
<< ntap >>
rect 1152 -44 1368 44
rect 1152 44 1368 132
rect 1152 132 1368 220
rect 1152 220 1368 308
rect 1152 308 1368 396
rect 1152 396 1368 484
rect 1152 484 1368 572
<< poly >>
rect 216 -36 936 36
rect 216 228 936 300
rect 216 492 936 564
rect 720 220 936 308
<< locali >>
rect 720 234 936 294
rect 1152 -44 1368 44
rect 1152 44 1368 132
rect 288 146 504 206
rect 288 146 504 206
rect 1152 132 1368 220
rect 720 234 936 294
rect 1152 220 1368 308
rect 1152 220 1368 308
rect 288 322 504 382
rect 288 322 504 382
rect 1152 308 1368 396
rect 1152 396 1368 484
rect 1152 484 1368 572
<< pcontact >>
rect 744 242 792 264
rect 744 264 792 286
rect 792 242 864 264
rect 792 264 864 286
rect 864 242 912 264
rect 864 264 912 286
<< ntapc >>
rect 1224 132 1296 220
rect 1224 308 1296 396
<< pdcontact >>
rect 312 154 360 176
rect 312 176 360 198
rect 360 154 432 176
rect 360 176 432 198
rect 432 154 480 176
rect 432 176 480 198
rect 312 330 360 352
rect 312 352 360 374
rect 360 330 432 352
rect 360 352 432 374
rect 432 330 480 352
rect 432 352 480 374
<< pmoslvt >>
rect 288 228 504 300
<< nwell >>
rect 0 -132 1440 660
<< labels >>
flabel locali s 720 234 936 294 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 288 146 504 206 0 FreeSans 400 0 0 0 S
port 3 nsew
flabel locali s 1152 220 1368 308 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 288 322 504 382 0 FreeSans 400 0 0 0 D
port 1 nsew
<< end >>
