magic
tech sky130A
magscale 1 2
timestamp 1658060514
<< checkpaint >>
rect 0 0 11760 4800
<< m1 >>
rect 2310 1810 2670 1870
rect 2400 530 2538 590
rect 2538 770 2760 830
rect 2538 530 2598 838
rect 360 2370 498 2430
rect 498 3090 1860 3150
rect 498 2370 558 3158
rect 1500 2050 1638 2110
rect 1638 2480 2400 2540
rect 1638 2050 1698 2552
rect 720 690 858 750
rect 858 1490 1860 1550
rect 858 690 918 1558
<< locali >>
rect 522 50 720 110
rect 522 370 720 430
rect 522 690 720 750
rect 522 1010 720 1070
rect 522 1330 720 1390
rect 522 1650 720 1710
rect 522 1970 720 2030
rect 522 2290 720 2350
rect 522 50 582 2350
rect 330 130 390 1150
rect 330 1410 390 2430
rect 720 210 858 270
rect 720 530 858 590
rect 720 850 858 910
rect 720 1170 858 1230
rect 858 210 918 1230
rect 720 1490 858 1550
rect 720 1810 858 1870
rect 720 2130 858 2190
rect 720 2450 858 2510
rect 858 1490 918 2510
<< m2 >>
rect 1500 1730 1638 1790
rect 1638 560 1860 620
rect 1638 560 1698 1798
rect 1134 2130 1860 2190
rect 360 770 1134 830
rect 1134 770 1194 2198
rect 2400 1330 2538 1390
rect 2538 -40 3482 20
rect 2538 -40 2598 1398
<< m3 >>
rect 3282 2680 7560 2740
rect 2762 1810 3282 1870
rect 3282 1810 3342 2740
rect 2310 0 2494 4800
rect 1770 0 1954 4800
use NCHDLR M1
transform 1 0 0 0 1 0
box 0 0 1140 320
use NCHDLR M2
transform 1 0 0 0 1 320
box 0 320 1140 640
use NCHDLR M3
transform 1 0 0 0 1 640
box 0 640 1140 960
use NCHDLR M4
transform 1 0 0 0 1 960
box 0 960 1140 1280
use NCHDLR M5
transform 1 0 0 0 1 1280
box 0 1280 1140 1600
use NCHDLR M6
transform 1 0 0 0 1 1600
box 0 1600 1140 1920
use NCHDLR M7
transform 1 0 0 0 1 1920
box 0 1920 1140 2240
use NCHDLR M8
transform 1 0 0 0 1 2240
box 0 2240 1140 2560
use TAPCELLB_CV XA5b
transform 1 0 1140 0 1 0
box 1140 0 3120 320
use IVX1_CV XA0
transform 1 0 1140 0 1 320
box 1140 320 3120 640
use TGPD_CV XA3
transform 1 0 1140 0 1 640
box 1140 640 3120 1600
use SARBSSWCTRL_CV XA4
transform 1 0 1140 0 1 1600
box 1140 1600 3120 2240
use TIEH_CV XA1
transform 1 0 1140 0 1 2240
box 1140 2240 3120 2560
use TAPCELLB_CV XA7
transform 1 0 1140 0 1 2560
box 1140 2560 3120 2880
use TIEL_CV XA2
transform 1 0 1140 0 1 2880
box 1140 2880 3120 3200
use TAPCELLB_CV XA5
transform 1 0 1140 0 1 3200
box 1140 3200 3120 3520
use CAP_BSSW5_CV XCAPB1
transform 1 0 3300 0 1 0
box 3300 0 11760 4800
use cut_M1M2_2x1 
transform 1 0 2310 0 1 1810
box 2310 1810 2494 1878
use cut_M2M4_2x1 
transform 1 0 2670 0 1 1810
box 2670 1810 2854 1878
use cut_M1M2_2x1 
transform 1 0 2310 0 1 530
box 2310 530 2494 598
use cut_M1M2_2x1 
transform 1 0 2670 0 1 770
box 2670 770 2854 838
use cut_M1M3_2x1 
transform 1 0 1410 0 1 1730
box 1410 1730 1594 1798
use cut_M1M3_2x1 
transform 1 0 1770 0 1 564
box 1770 564 1954 632
use cut_M1M2_2x1 
transform 1 0 270 0 1 2370
box 270 2370 454 2438
use cut_M1M2_2x1 
transform 1 0 1770 0 1 3090
box 1770 3090 1954 3158
use cut_M1M2_2x1 
transform 1 0 1410 0 1 2050
box 1410 2050 1594 2118
use cut_M1M2_2x1 
transform 1 0 2310 0 1 2484
box 2310 2484 2494 2552
use cut_M1M2_2x1 
transform 1 0 630 0 1 690
box 630 690 814 758
use cut_M1M2_2x1 
transform 1 0 1770 0 1 1490
box 1770 1490 1954 1558
use cut_M1M3_2x1 
transform 1 0 1766 0 1 2130
box 1766 2130 1950 2198
use cut_M1M3_2x1 
transform 1 0 266 0 1 770
box 266 770 450 838
use cut_M1M3_2x1 
transform 1 0 2310 0 1 1330
box 2310 1330 2494 1398
use cut_M3M4_2x1 
transform 1 0 3390 0 1 -40
box 3390 -40 3574 28
use cut_M1M4_2x1 
transform 1 0 626 0 1 46
box 626 46 810 114
use cut_M2M4_2x1 
transform 1 0 1214 0 1 3086
box 1214 3086 1398 3154
<< labels >>
flabel m3 s 626 46 810 114 0 FreeSans 400 0 0 0 VI
port 1 nsew
flabel m3 s 1214 3086 1398 3154 0 FreeSans 400 0 0 0 TIE_L
port 2 nsew
flabel locali s 1410 450 1590 510 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel locali s 2670 770 2850 830 0 FreeSans 400 0 0 0 CKN
port 4 nsew
flabel locali s 630 1170 810 1230 0 FreeSans 400 0 0 0 VO1
port 5 nsew
flabel locali s 630 2450 810 2510 0 FreeSans 400 0 0 0 VO2
port 6 nsew
flabel m3 s 2310 0 2494 4800 0 FreeSans 400 0 0 0 AVDD
port 7 nsew
flabel m3 s 1770 0 1954 4800 0 FreeSans 400 0 0 0 AVSS
port 8 nsew
<< end >>
