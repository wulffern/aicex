magic
tech sky130A
magscale 1 2
timestamp 1660740729
<< checkpaint >>
rect -640 -640 1288 3500
<< locali >>
rect -640 -640 1288 -528
rect -640 -640 1288 -528
rect -640 -640 -528 3500
rect -640 3388 1288 3500
rect 1176 -640 1288 3500
rect -640 -640 1288 -528
rect 378 2750 702 2970
rect -54 2750 270 2970
<< ptapc >>
rect -636 -640 -556 -560
rect -556 -640 -476 -560
rect -476 -640 -396 -560
rect -396 -640 -316 -560
rect -316 -640 -236 -560
rect -236 -640 -156 -560
rect -156 -640 -76 -560
rect -76 -640 4 -560
rect 4 -640 84 -560
rect 84 -640 164 -560
rect 164 -640 244 -560
rect 244 -640 324 -560
rect 324 -640 404 -560
rect 404 -640 484 -560
rect 484 -640 564 -560
rect 564 -640 644 -560
rect 644 -640 724 -560
rect 724 -640 804 -560
rect 804 -640 884 -560
rect 884 -640 964 -560
rect 964 -640 1044 -560
rect 1044 -640 1124 -560
rect 1124 -640 1204 -560
rect 1204 -640 1284 -560
rect -640 -610 -560 -530
rect -640 -530 -560 -450
rect -640 -450 -560 -370
rect -640 -370 -560 -290
rect -640 -290 -560 -210
rect -640 -210 -560 -130
rect -640 -130 -560 -50
rect -640 -50 -560 30
rect -640 30 -560 110
rect -640 110 -560 190
rect -640 190 -560 270
rect -640 270 -560 350
rect -640 350 -560 430
rect -640 430 -560 510
rect -640 510 -560 590
rect -640 590 -560 670
rect -640 670 -560 750
rect -640 750 -560 830
rect -640 830 -560 910
rect -640 910 -560 990
rect -640 990 -560 1070
rect -640 1070 -560 1150
rect -640 1150 -560 1230
rect -640 1230 -560 1310
rect -640 1310 -560 1390
rect -640 1390 -560 1470
rect -640 1470 -560 1550
rect -640 1550 -560 1630
rect -640 1630 -560 1710
rect -640 1710 -560 1790
rect -640 1790 -560 1870
rect -640 1870 -560 1950
rect -640 1950 -560 2030
rect -640 2030 -560 2110
rect -640 2110 -560 2190
rect -640 2190 -560 2270
rect -640 2270 -560 2350
rect -640 2350 -560 2430
rect -640 2430 -560 2510
rect -640 2510 -560 2590
rect -640 2590 -560 2670
rect -640 2670 -560 2750
rect -640 2750 -560 2830
rect -640 2830 -560 2910
rect -640 2910 -560 2990
rect -640 2990 -560 3070
rect -640 3070 -560 3150
rect -640 3150 -560 3230
rect -640 3230 -560 3310
rect -640 3310 -560 3390
rect -640 3390 -560 3470
rect -636 3388 -556 3468
rect -556 3388 -476 3468
rect -476 3388 -396 3468
rect -396 3388 -316 3468
rect -316 3388 -236 3468
rect -236 3388 -156 3468
rect -156 3388 -76 3468
rect -76 3388 4 3468
rect 4 3388 84 3468
rect 84 3388 164 3468
rect 164 3388 244 3468
rect 244 3388 324 3468
rect 324 3388 404 3468
rect 404 3388 484 3468
rect 484 3388 564 3468
rect 564 3388 644 3468
rect 644 3388 724 3468
rect 724 3388 804 3468
rect 804 3388 884 3468
rect 884 3388 964 3468
rect 964 3388 1044 3468
rect 1044 3388 1124 3468
rect 1124 3388 1204 3468
rect 1204 3388 1284 3468
rect 1176 -610 1256 -530
rect 1176 -530 1256 -450
rect 1176 -450 1256 -370
rect 1176 -370 1256 -290
rect 1176 -290 1256 -210
rect 1176 -210 1256 -130
rect 1176 -130 1256 -50
rect 1176 -50 1256 30
rect 1176 30 1256 110
rect 1176 110 1256 190
rect 1176 190 1256 270
rect 1176 270 1256 350
rect 1176 350 1256 430
rect 1176 430 1256 510
rect 1176 510 1256 590
rect 1176 590 1256 670
rect 1176 670 1256 750
rect 1176 750 1256 830
rect 1176 830 1256 910
rect 1176 910 1256 990
rect 1176 990 1256 1070
rect 1176 1070 1256 1150
rect 1176 1150 1256 1230
rect 1176 1230 1256 1310
rect 1176 1310 1256 1390
rect 1176 1390 1256 1470
rect 1176 1470 1256 1550
rect 1176 1550 1256 1630
rect 1176 1630 1256 1710
rect 1176 1710 1256 1790
rect 1176 1790 1256 1870
rect 1176 1870 1256 1950
rect 1176 1950 1256 2030
rect 1176 2030 1256 2110
rect 1176 2110 1256 2190
rect 1176 2190 1256 2270
rect 1176 2270 1256 2350
rect 1176 2350 1256 2430
rect 1176 2430 1256 2510
rect 1176 2510 1256 2590
rect 1176 2590 1256 2670
rect 1176 2670 1256 2750
rect 1176 2750 1256 2830
rect 1176 2830 1256 2910
rect 1176 2910 1256 2990
rect 1176 2990 1256 3070
rect 1176 3070 1256 3150
rect 1176 3150 1256 3230
rect 1176 3230 1256 3310
rect 1176 3310 1256 3390
rect 1176 3390 1256 3470
<< ptap >>
rect -640 -640 1288 -528
rect -640 -640 -528 3500
rect -640 3388 1288 3500
rect 1176 -640 1288 3500
use SUNTR_RES12 XA1
transform 1 0 0 0 1 0
box 0 0 648 2860
<< labels >>
flabel locali s -640 -640 1288 -528 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 378 2750 702 2970 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s -54 2750 270 2970 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
