magic
tech sky130A
magscale 1 2
timestamp 1660114332
<< checkpaint >>
rect 0 0 1260 528
<< locali >>
rect 864 58 1032 118
rect 864 410 1032 470
rect 1032 58 1092 470
rect 402 146 462 382
rect -108 132 108 220
rect 756 234 972 294
rect 324 146 540 206
rect 756 58 972 118
use SUNTR_NCHDL M0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_NCHDL M1
transform 1 0 0 0 1 176
box 0 176 1260 528
<< labels >>
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 756 234 972 294 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 756 58 972 118 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
