magic
tech sky130A
magscale 1 2
timestamp 1660085871
<< checkpaint >>
rect -108 -896 2520 2992
<< m2 >>
rect 0 -448 2520 -144
rect 0 -448 2520 -144
rect 0 -896 2520 -592
rect 0 -896 2520 -592
<< m3 >>
rect 748 -448 964 704
rect 1540 -896 1756 704
<< locali >>
rect 432 1026 600 1086
rect 600 586 864 646
rect 600 586 660 1086
rect 636 1174 816 1234
rect 636 2874 864 2934
rect 432 1378 636 1438
rect 636 1174 696 2934
rect 756 1114 864 1174
rect -108 352 108 1452
rect 756 1114 972 1174
rect 324 498 540 558
<< m1 >>
rect 864 938 1032 998
rect 864 1290 1032 1350
rect 856 352 1032 412
rect 1032 352 1092 1358
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV xa00
transform 1 0 0 0 1 0
box 0 0 2520 352
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV xa10
transform 1 0 0 0 1 352
box 0 352 2520 704
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa20
transform 1 0 0 0 1 880
box 0 880 1260 1232
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa30
transform 1 0 0 0 1 1232
box 0 1232 1260 2992
use cut_M3M4_2x1 
transform 1 0 756 0 1 -448
box 756 -448 956 -372
use cut_M3M4_2x1 
transform 1 0 1548 0 1 -896
box 1548 -896 1748 -820
use cut_M1M2_2x1 
transform 1 0 788 0 1 938
box 788 938 972 1006
use cut_M1M2_2x1 
transform 1 0 788 0 1 1290
box 788 1290 972 1358
use cut_M1M4_1x2 
transform 1 0 -38 0 1 352
box -38 352 38 552
<< labels >>
flabel m2 s 0 -448 2520 -144 0 FreeSans 400 0 0 0 AVSS
port 4 nsew
flabel m2 s 0 -896 2520 -592 0 FreeSans 400 0 0 0 AVDD
port 2 nsew
flabel locali s 756 1114 972 1174 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
<< end >>
