magic
tech sky130A
magscale 1 2
timestamp 1657978845
<< checkpaint >>
rect 0 0 2320 2240
<< poly >>
rect 280 2062 2040 2098
rect 280 142 2040 178
<< locali >>
rect 1890 1410 1950 2110
rect 370 450 430 1790
rect 800 530 968 590
rect 800 1170 968 1230
rect 800 1810 968 1870
rect 968 530 1520 590
rect 968 530 1028 1870
rect 572 210 800 270
rect 572 850 800 910
rect 572 1490 800 1550
rect 572 210 632 1550
rect 800 210 968 270
rect 968 50 1520 110
rect 968 50 1028 270
rect 1292 1170 1520 1230
rect 1292 1810 1520 1870
rect 800 2130 1292 2190
rect 1292 1170 1352 2190
rect 1920 130 2088 190
rect 1920 450 2088 510
rect 1920 1090 2088 1150
rect 2088 130 2148 1150
rect 770 210 830 430
rect 770 530 830 750
rect 770 850 830 1070
rect 770 1170 830 1390
rect 770 1490 830 1710
rect 770 1810 830 2030
rect 1490 210 1550 430
rect 1490 530 1550 750
rect 1490 850 1550 1070
rect 1490 1170 1550 1390
rect 1490 1490 1550 1710
rect 1490 1810 1550 2030
<< m3 >>
rect 1520 850 1688 910
rect 1688 770 1920 830
rect 1688 770 1748 918
rect 1400 0 1600 2240
rect 680 0 880 2240
use NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1160 320
use NCHDL MN1
transform 1 0 0 0 1 320
box 0 320 1160 640
use NCHDL MN2
transform 1 0 0 0 1 640
box 0 640 1160 960
use NCHDL MN3
transform 1 0 0 0 1 960
box 0 960 1160 1280
use NCHDL MN4
transform 1 0 0 0 1 1280
box 0 1280 1160 1600
use NCHDL MN5
transform 1 0 0 0 1 1600
box 0 1600 1160 1920
use NCHDL MN6
transform 1 0 0 0 1 1920
box 0 1920 1160 2240
use PCHDL MP0
transform 1 0 1160 0 1 0
box 1160 0 2320 320
use PCHDL MP1
transform 1 0 1160 0 1 320
box 1160 320 2320 640
use PCHDL MP2
transform 1 0 1160 0 1 640
box 1160 640 2320 960
use PCHDL MP3
transform 1 0 1160 0 1 960
box 1160 960 2320 1280
use PCHDL MP4
transform 1 0 1160 0 1 1280
box 1160 1280 2320 1600
use PCHDL MP5
transform 1 0 1160 0 1 1600
box 1160 1600 2320 1920
use PCHDL MP6
transform 1 0 1160 0 1 1920
box 1160 1920 2320 2240
use cut_M1M4_2x1 
transform 1 0 1400 0 1 850
box 1400 850 1600 918
use cut_M1M4_2x1 
transform 1 0 1800 0 1 770
box 1800 770 2000 838
use cut_M1M4_2x1 
transform 1 0 1400 0 1 210
box 1400 210 1600 278
use cut_M1M4_2x1 
transform 1 0 1400 0 1 370
box 1400 370 1600 438
use cut_M1M4_2x1 
transform 1 0 1400 0 1 850
box 1400 850 1600 918
use cut_M1M4_2x1 
transform 1 0 1400 0 1 1010
box 1400 1010 1600 1078
use cut_M1M4_2x1 
transform 1 0 1400 0 1 1490
box 1400 1490 1600 1558
use cut_M1M4_2x1 
transform 1 0 1400 0 1 1650
box 1400 1650 1600 1718
use cut_M1M4_2x1 
transform 1 0 1400 0 1 2130
box 1400 2130 1600 2198
use cut_M1M4_2x1 
transform 1 0 680 0 1 50
box 680 50 880 118
<< labels >>
flabel locali s 2200 120 2440 200 0 FreeSans 400 0 0 0 BULKP
port 1 nsew
flabel locali s -120 120 120 200 0 FreeSans 400 0 0 0 BULKN
port 2 nsew
flabel locali s 680 1490 920 1550 0 FreeSans 400 0 0 0 N1
port 3 nsew
flabel locali s 680 1810 920 1870 0 FreeSans 400 0 0 0 N2
port 4 nsew
flabel locali s 280 450 520 510 0 FreeSans 400 0 0 0 CI
port 5 nsew
flabel locali s 280 130 520 190 0 FreeSans 400 0 0 0 CK
port 6 nsew
flabel locali s 680 2130 920 2190 0 FreeSans 400 0 0 0 CO
port 7 nsew
flabel locali s 280 2050 520 2110 0 FreeSans 400 0 0 0 VMR
port 8 nsew
flabel m3 s 1400 0 1600 2240 0 FreeSans 400 0 0 0 AVDD
port 9 nsew
flabel m3 s 680 0 880 2240 0 FreeSans 400 0 0 0 AVSS
port 10 nsew
<< end >>
