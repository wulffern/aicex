magic
tech sky130A
magscale 1 2
timestamp 1658699483
<< checkpaint >>
rect 0 30 9504 2870
<< m3 >>
rect 328 0 404 2900
rect 328 0 404 2900
rect 468 140 544 2760
rect 608 0 684 2900
rect 748 140 824 2760
rect 888 0 964 2900
rect 1028 140 1104 2760
rect 1168 0 1244 2900
rect 1308 140 1384 2760
rect 1448 0 1524 2900
rect 1588 140 1664 2760
rect 1728 0 1804 2900
rect 1868 140 1944 2760
rect 2008 0 2084 2900
rect 2148 140 2224 2760
rect 2288 0 2364 2900
rect 2428 140 2504 2760
rect 2568 0 2644 2900
rect 2708 140 2784 2760
rect 2848 0 2924 2900
rect 2988 140 3064 2760
rect 3128 0 3204 2900
rect 3268 140 3344 2760
rect 3408 0 3484 2900
rect 3548 140 3624 2760
rect 3688 0 3764 2900
rect 3828 140 3904 2760
rect 3968 0 4044 2900
rect 4108 140 4184 2760
rect 4248 0 4324 2900
rect 4388 140 4464 2760
rect 4528 0 4604 2900
rect 4668 140 4744 2760
rect 4808 0 4884 2900
rect 4948 140 5024 2760
rect 5088 0 5164 2900
rect 5228 140 5304 2760
rect 5368 0 5444 2900
rect 5508 140 5584 2760
rect 5648 0 5724 2900
rect 5788 140 5864 2760
rect 5928 0 6004 2900
rect 6068 140 6144 2760
rect 6208 0 6284 2900
rect 6348 140 6424 2760
rect 6488 0 6564 2900
rect 6628 140 6704 2760
rect 6768 0 6844 2900
rect 6908 140 6984 2760
rect 7048 0 7124 2900
rect 7188 140 7264 2760
rect 7328 0 7404 2900
rect 7468 140 7544 2760
rect 7608 0 7684 2900
rect 7748 140 7824 2760
rect 7888 0 7964 2900
rect 8028 140 8104 2760
rect 8168 0 8244 2900
rect 8308 140 8384 2760
rect 8448 0 8524 2900
rect 8588 140 8664 2760
rect 8728 0 8804 2900
rect 8868 140 8944 2760
rect 9008 0 9084 2900
rect 9148 140 9224 2760
rect 9428 0 9504 2900
rect 9288 0 9364 2900
rect 328 0 9288 76
rect 328 2824 9288 2900
<< m1 >>
rect 328 0 9428 76
rect 2428 400 2504 2900
rect 7188 0 7264 2500
rect 2708 0 2784 1048
rect 2708 1368 2784 2900
rect 6908 0 6984 1048
rect 6908 1368 6984 2900
rect 2148 0 2224 2016
rect 2148 2336 2224 2900
rect 2988 0 3064 2016
rect 2988 2336 3064 2900
rect 6628 0 6704 2016
rect 6628 2336 6704 2900
rect 7468 0 7544 2016
rect 7468 2336 7544 2900
rect 1588 0 1664 1532
rect 1588 1852 1664 2900
rect 1868 0 1944 1532
rect 1868 1852 1944 2900
rect 3268 0 3344 1532
rect 3268 1852 3344 2900
rect 3548 0 3624 1532
rect 3548 1852 3624 2900
rect 6068 0 6144 1532
rect 6068 1852 6144 2900
rect 6348 0 6424 1532
rect 6348 1852 6424 2900
rect 7748 0 7824 1532
rect 7748 1852 7824 2900
rect 8028 0 8104 1532
rect 8028 1852 8104 2900
rect 468 0 544 564
rect 468 884 544 2900
rect 748 0 824 564
rect 748 884 824 2900
rect 1028 0 1104 564
rect 1028 884 1104 2900
rect 1308 0 1384 564
rect 1308 884 1384 2900
rect 3828 0 3904 564
rect 3828 884 3904 2900
rect 4108 0 4184 564
rect 4108 884 4184 2900
rect 4388 0 4464 564
rect 4388 884 4464 2900
rect 4668 0 4744 564
rect 4668 884 4744 2900
rect 4948 0 5024 564
rect 4948 884 5024 2900
rect 5228 0 5304 564
rect 5228 884 5304 2900
rect 5508 0 5584 564
rect 5508 884 5584 2900
rect 5788 0 5864 564
rect 5788 884 5864 2900
rect 8308 0 8384 564
rect 8308 884 8384 2900
rect 8588 0 8664 564
rect 8588 884 8664 2900
rect 8868 0 8944 564
rect 8868 884 8944 2900
rect 9148 0 9224 564
rect 9148 884 9224 2900
rect 328 0 404 2824
rect 608 0 684 2824
rect 888 0 964 2824
rect 1168 0 1244 2824
rect 1448 0 1524 2824
rect 1728 0 1804 2824
rect 2008 0 2084 2824
rect 2288 0 2364 2824
rect 2568 0 2644 2824
rect 2848 0 2924 2824
rect 3128 0 3204 2824
rect 3408 0 3484 2824
rect 3688 0 3764 2824
rect 3968 0 4044 2824
rect 4248 0 4324 2824
rect 4528 0 4604 2824
rect 4808 0 4884 2824
rect 5088 0 5164 2824
rect 5368 0 5444 2824
rect 5648 0 5724 2824
rect 5928 0 6004 2824
rect 6208 0 6284 2824
rect 6488 0 6564 2824
rect 6768 0 6844 2824
rect 7048 0 7124 2824
rect 7328 0 7404 2824
rect 7608 0 7684 2824
rect 7888 0 7964 2824
rect 8168 0 8244 2824
rect 8448 0 8524 2824
rect 8728 0 8804 2824
rect 9008 0 9084 2824
rect 9428 0 9504 2900
rect 9288 0 9364 2900
rect 328 0 9428 76
rect 328 2824 9428 2900
<< locali >>
rect 0 202 200 278
rect 0 2622 200 2698
rect 0 1170 200 1246
rect 0 2138 200 2214
rect 0 1654 200 1730
rect 0 686 200 762
rect 320 686 9288 762
rect 320 202 9288 278
rect 320 2622 9288 2698
rect 320 1170 9288 1246
rect 320 2138 9288 2214
rect 320 1654 9288 1730
<< m4 >>
rect 188 0 264 2900
rect 468 0 544 2900
rect 748 0 824 2900
rect 1028 0 1104 2900
rect 1308 0 1384 2900
rect 1588 0 1664 2900
rect 1868 0 1944 2900
rect 2148 0 2224 2900
rect 2428 0 2504 2900
rect 2708 0 2784 2900
rect 2988 0 3064 2900
rect 3268 0 3344 2900
rect 3548 0 3624 2900
rect 3828 0 3904 2900
rect 4108 0 4184 2900
rect 4388 0 4464 2900
rect 4668 0 4744 2900
rect 4948 0 5024 2900
rect 5228 0 5304 2900
rect 5508 0 5584 2900
rect 5788 0 5864 2900
rect 6068 0 6144 2900
rect 6348 0 6424 2900
rect 6628 0 6704 2900
rect 6908 0 6984 2900
rect 7188 0 7264 2900
rect 7468 0 7544 2900
rect 7748 0 7824 2900
rect 8028 0 8104 2900
rect 8308 0 8384 2900
rect 8588 0 8664 2900
rect 8868 0 8944 2900
rect 9148 0 9224 2900
rect 9428 0 9504 2900
rect 188 0 9428 76
rect 188 2824 9428 2900
<< m2 >>
rect 9428 0 9504 2900
use RM1 XRES1A
transform 1 0 200 0 1 202
box 200 202 320 202
use RM1 XRES1B
transform 1 0 200 0 1 2622
box 200 2622 320 2622
use RM1 XRES2
transform 1 0 200 0 1 1170
box 200 1170 320 1170
use RM1 XRES4
transform 1 0 200 0 1 2138
box 200 2138 320 2138
use RM1 XRES8
transform 1 0 200 0 1 1654
box 200 1654 320 1654
use RM1 XRES16
transform 1 0 200 0 1 686
box 200 686 320 686
use cut_M2M5_1x2 
transform 1 0 9428 0 1 1250
box 9428 1250 9504 1450
use cut_M1M4_1x2 
transform 1 0 2428 0 1 140
box 2428 140 2504 340
use cut_M1M4_1x2 
transform 1 0 7188 0 1 2560
box 7188 2560 7264 2760
use cut_M1M4_1x2 
transform 1 0 2708 0 1 1108
box 2708 1108 2784 1308
use cut_M1M4_1x2 
transform 1 0 6908 0 1 1108
box 6908 1108 6984 1308
use cut_M1M4_1x2 
transform 1 0 2148 0 1 2076
box 2148 2076 2224 2276
use cut_M1M4_1x2 
transform 1 0 2988 0 1 2076
box 2988 2076 3064 2276
use cut_M1M4_1x2 
transform 1 0 6628 0 1 2076
box 6628 2076 6704 2276
use cut_M1M4_1x2 
transform 1 0 7468 0 1 2076
box 7468 2076 7544 2276
use cut_M1M4_1x2 
transform 1 0 1588 0 1 1592
box 1588 1592 1664 1792
use cut_M1M4_1x2 
transform 1 0 1868 0 1 1592
box 1868 1592 1944 1792
use cut_M1M4_1x2 
transform 1 0 3268 0 1 1592
box 3268 1592 3344 1792
use cut_M1M4_1x2 
transform 1 0 3548 0 1 1592
box 3548 1592 3624 1792
use cut_M1M4_1x2 
transform 1 0 6068 0 1 1592
box 6068 1592 6144 1792
use cut_M1M4_1x2 
transform 1 0 6348 0 1 1592
box 6348 1592 6424 1792
use cut_M1M4_1x2 
transform 1 0 7748 0 1 1592
box 7748 1592 7824 1792
use cut_M1M4_1x2 
transform 1 0 8028 0 1 1592
box 8028 1592 8104 1792
use cut_M1M4_1x2 
transform 1 0 468 0 1 624
box 468 624 544 824
use cut_M1M4_1x2 
transform 1 0 748 0 1 624
box 748 624 824 824
use cut_M1M4_1x2 
transform 1 0 1028 0 1 624
box 1028 624 1104 824
use cut_M1M4_1x2 
transform 1 0 1308 0 1 624
box 1308 624 1384 824
use cut_M1M4_1x2 
transform 1 0 3828 0 1 624
box 3828 624 3904 824
use cut_M1M4_1x2 
transform 1 0 4108 0 1 624
box 4108 624 4184 824
use cut_M1M4_1x2 
transform 1 0 4388 0 1 624
box 4388 624 4464 824
use cut_M1M4_1x2 
transform 1 0 4668 0 1 624
box 4668 624 4744 824
use cut_M1M4_1x2 
transform 1 0 4948 0 1 624
box 4948 624 5024 824
use cut_M1M4_1x2 
transform 1 0 5228 0 1 624
box 5228 624 5304 824
use cut_M1M4_1x2 
transform 1 0 5508 0 1 624
box 5508 624 5584 824
use cut_M1M4_1x2 
transform 1 0 5788 0 1 624
box 5788 624 5864 824
use cut_M1M4_1x2 
transform 1 0 8308 0 1 624
box 8308 624 8384 824
use cut_M1M4_1x2 
transform 1 0 8588 0 1 624
box 8588 624 8664 824
use cut_M1M4_1x2 
transform 1 0 8868 0 1 624
box 8868 624 8944 824
use cut_M1M4_1x2 
transform 1 0 9148 0 1 624
box 9148 624 9224 824
<< labels >>
flabel m3 s 328 0 404 2900 0 FreeSans 400 0 0 0 CTOP
port 7 nsew
flabel m1 s 328 0 9428 76 0 FreeSans 400 0 0 0 AVSS
port 8 nsew
flabel locali s 0 202 200 278 0 FreeSans 400 0 0 0 C1A
port 1 nsew
flabel locali s 0 2622 200 2698 0 FreeSans 400 0 0 0 C1B
port 2 nsew
flabel locali s 0 1170 200 1246 0 FreeSans 400 0 0 0 C2
port 3 nsew
flabel locali s 0 2138 200 2214 0 FreeSans 400 0 0 0 C4
port 4 nsew
flabel locali s 0 1654 200 1730 0 FreeSans 400 0 0 0 C8
port 5 nsew
flabel locali s 0 686 200 762 0 FreeSans 400 0 0 0 C16
port 6 nsew
<< end >>
