magic
tech sky130A
magscale 1 2
timestamp 1658072521
<< checkpaint >>
rect -1736 -1560 24904 39226
<< m3 >>
rect 8580 17456 23334 17524
rect 8580 17836 23334 17904
rect 21634 18176 21702 25396
rect 21878 18176 21946 32436
rect 4834 18284 4902 28592
rect 5550 18474 5618 28592
rect 9034 18664 9102 28592
rect 1350 18854 1418 28592
rect 1350 18854 1418 28592
rect 12738 19044 12806 28614
rect 12738 19044 12806 28614
rect 16938 19234 17006 28614
rect 16938 19234 17006 28614
rect 10362 19424 10430 28614
rect 10362 19424 10430 28614
rect 14562 19614 14630 28614
rect 14562 19614 14630 28614
rect 1962 19804 2030 28614
rect 6162 19994 6230 28614
rect 6162 19994 6230 28614
rect 4338 20184 4406 28614
rect 4338 20184 4406 28614
rect 8538 20374 8606 28614
rect 8538 20374 8606 28614
rect 2098 20564 2166 29894
rect 8402 20754 8470 29894
rect 6298 20944 6366 29894
rect 4202 21134 4270 29894
rect 10634 21324 10702 31174
rect 12466 21514 12534 31174
rect 14834 21704 14902 31174
rect 8266 21894 8334 31174
rect 4066 22084 4134 31174
rect 2234 22274 2302 31174
rect 16666 22464 16734 31174
rect 6434 22654 6502 31174
rect 1714 23346 1898 38026
rect 4470 23346 4654 38026
rect 5914 23346 6098 38026
rect 8670 23346 8854 38026
rect 10114 23346 10298 38026
rect 12870 23346 13054 38026
rect 14314 23346 14498 38026
rect 17070 23346 17254 38026
rect 18514 23346 18698 38026
rect 21270 23346 21454 38026
rect 9570 -600 9754 4800
rect 13414 -600 13598 4800
rect 2374 23346 2558 38626
rect 3810 23346 3994 38626
rect 6574 23346 6758 38626
rect 8010 23346 8194 38626
rect 10774 23346 10958 38626
rect 12210 23346 12394 38626
rect 14974 23346 15158 38626
rect 16410 23346 16594 38626
rect 19174 23346 19358 38626
rect 20610 23346 20794 38626
rect 8910 -1200 9094 4800
rect 14074 -1200 14258 4800
rect 2854 27716 3038 39226
rect 3330 27716 3514 39226
rect 7054 27716 7238 39226
rect 7530 27716 7714 39226
rect 11254 27716 11438 39226
rect 11730 27716 11914 39226
rect 15454 27716 15638 39226
rect 15930 27716 16114 39226
rect 19654 27716 19838 39226
rect 10184 -1560 10252 3154
rect 12916 -1560 12984 3154
rect 10642 1170 10864 1238
rect 8614 4990 10642 5058
rect 12304 1170 12458 1238
rect 12458 4990 14534 5058
rect 10864 1170 11018 1238
rect 11018 2450 12304 2518
rect 11018 1170 11086 2518
rect 10774 46 10958 114
rect 12210 46 12394 114
rect 18762 28614 18830 28798
<< m2 >>
rect 14500 16954 14568 17524
rect 8580 16954 8648 17904
rect 4834 18216 13624 18284
rect 5550 18406 13248 18474
rect 9034 18596 12872 18664
rect 1350 18786 14000 18854
rect 10848 18976 12806 19044
rect 11224 19166 17006 19234
rect 10362 19356 10728 19424
rect 11036 19546 14630 19614
rect 1962 19736 9224 19804
rect 6162 19926 9976 19994
rect 4338 20116 9600 20184
rect 8538 20306 10352 20374
rect 2098 20496 9412 20564
rect 8402 20686 10540 20754
rect 6298 20876 10164 20944
rect 4202 21066 9788 21134
rect 10634 21256 12496 21324
rect 12240 21446 12534 21514
rect 12052 21636 14902 21704
rect 8266 21826 12684 21894
rect 4066 22016 13436 22084
rect 2234 22206 13812 22274
rect 11864 22396 16734 22464
rect 6434 22586 13060 22654
rect 2374 36066 2682 36134
rect 2682 35504 4834 35572
rect 4766 35504 4834 35696
rect 2682 35504 2750 36138
rect 6574 36066 6882 36134
rect 6882 35504 9034 35572
rect 8966 35504 9034 35696
rect 6882 35504 6950 36138
rect 10774 36066 11082 36134
rect 11082 35504 13234 35572
rect 13166 35504 13234 35696
rect 11082 35504 11150 36138
rect 14974 36066 15282 36134
rect 15282 35504 17434 35572
rect 17366 35504 17434 35696
rect 15282 35504 15350 36138
rect 1354 32624 18334 32692
rect 1286 32624 1354 32816
rect 4766 32624 4834 32816
rect 5486 32624 5554 32816
rect 8966 32624 9034 32816
rect 9686 32624 9754 32816
rect 13166 32624 13234 32816
rect 13886 32624 13954 32816
rect 17366 32624 17434 32816
rect 18086 32624 18154 32816
rect 2370 24032 2682 24100
rect 2682 23660 4834 23728
rect 4766 23660 4834 23860
rect 2682 23660 2750 24100
rect 6570 24032 6882 24100
rect 6882 23660 9034 23728
rect 8966 23660 9034 23860
rect 6882 23660 6950 24100
rect 10770 24032 11082 24100
rect 11082 23660 13234 23728
rect 13166 23660 13234 23860
rect 11082 23660 11150 24100
rect 14970 24032 15282 24100
rect 15282 23660 17434 23728
rect 17366 23660 17434 23860
rect 15282 23660 15350 24100
rect 19170 24032 19482 24100
rect 19482 24032 19550 24100
rect 3814 24032 4126 24100
rect 4126 24032 4194 24164
rect 4126 24164 5550 24232
rect 5482 23792 5550 24232
rect 8014 24032 8326 24100
rect 8326 24032 8394 24164
rect 8326 24164 9750 24232
rect 9682 23792 9750 24232
rect 12214 24032 12526 24100
rect 12526 24032 12594 24164
rect 12526 24164 13950 24232
rect 13882 23792 13950 24232
rect 16414 24032 16726 24100
rect 16726 24032 16794 24164
rect 16726 24164 18150 24232
rect 18082 23792 18150 24232
rect 1350 25748 18334 25816
rect 1282 25392 1350 25816
rect 4766 25392 4834 25816
rect 5482 25392 5550 25816
rect 8966 25392 9034 25816
rect 9682 25392 9750 25816
rect 13166 25392 13234 25816
rect 13882 25392 13950 25816
rect 17366 25392 17434 25816
rect 18082 25392 18150 25816
rect 1354 26000 18334 26068
rect 1286 26000 1354 26416
rect 4766 26000 4834 26416
rect 5486 26000 5554 26416
rect 8966 26000 9034 26416
rect 9686 26000 9754 26416
rect 13166 26000 13234 26416
rect 13886 26000 13954 26416
rect 17366 26000 17434 26416
rect 18086 26000 18154 26416
rect 2734 26996 1534 27056
rect 2734 26996 2914 27056
rect 2734 26996 3634 27056
rect 2734 26996 7114 27056
rect 2734 26996 7834 27056
rect 2734 26996 11314 27056
rect 2734 26996 12034 27056
rect 2734 26996 15514 27056
rect 2734 26996 16234 27056
rect 2734 26996 19714 27056
rect 21142 28386 21364 28454
rect 18266 25460 21142 25528
rect 21142 25460 21210 28458
rect 18242 25392 18334 25460
rect 20482 29666 20704 29734
rect 18266 26424 20482 26492
rect 20482 26424 20550 29738
rect 18244 26356 18334 26424
rect 20344 36276 20498 36344
rect 18244 33396 20498 33464
rect 20498 33396 20566 36344
rect 20122 36916 20344 36984
rect 19264 36066 20122 36134
rect 20122 36066 20190 36984
rect 10864 2450 11018 2518
rect 11018 1170 12304 1238
rect 11018 1170 11086 2518
rect 1354 26996 2914 27056
<< m4 >>
rect 21634 17836 21702 18176
rect 21878 17456 21946 18176
rect 10642 1170 10710 5058
rect 12458 1170 12526 5058
<< m1 >>
rect 13556 16894 13624 18216
rect 13180 16894 13248 18406
rect 12804 16894 12872 18596
rect 13932 16894 14000 18786
rect 10848 16894 10916 18976
rect 11224 16894 11292 19166
rect 10660 16894 10728 19356
rect 11036 16894 11104 19546
rect 9156 16894 9224 19736
rect 9908 16894 9976 19926
rect 9532 16894 9600 20116
rect 10284 16894 10352 20306
rect 9344 16894 9412 20496
rect 10472 16894 10540 20686
rect 10096 16894 10164 20876
rect 9720 16894 9788 21066
rect 12428 16894 12496 21256
rect 12240 16894 12308 21446
rect 12052 16894 12120 21636
rect 12616 16894 12684 21826
rect 13368 16894 13436 22016
rect 13744 16894 13812 22206
rect 11864 16894 11932 22396
rect 12992 16894 13060 22586
rect 9994 -1380 10054 510
rect 13114 -1380 13174 510
rect 1354 35636 -1676 35696
rect 3814 36036 4122 36096
rect 4122 35512 5554 35572
rect 5494 35512 5554 35696
rect 4122 35512 4182 36104
rect 8014 36036 8322 36096
rect 8322 35512 9754 35572
rect 9694 35512 9754 35696
rect 8322 35512 8382 36104
rect 12214 36036 12522 36096
rect 12522 35512 13954 35572
rect 13894 35512 13954 35696
rect 12522 35512 12582 36104
rect 16414 36036 16722 36096
rect 16722 35512 18154 35572
rect 18094 35512 18154 35696
rect 16722 35512 16782 36104
rect 20130 36596 20344 36656
rect 18604 34116 20130 34176
rect 20130 34116 20190 36664
rect -956 4990 68 5050
rect -956 6478 68 6538
rect -956 7966 68 8026
rect -956 9454 68 9514
rect -956 10942 68 11002
rect -956 12430 68 12490
rect -956 13918 68 13978
rect -956 15406 68 15466
rect 23080 4990 24124 5050
rect 23080 6478 24124 6538
rect 23080 7966 24124 8026
rect 23080 9454 24124 9514
rect 23080 10942 24124 11002
rect 23080 12430 24124 12490
rect 23080 13918 24124 13978
rect 23080 15406 24124 15466
<< locali >>
rect 23940 -600 24124 38026
rect -956 -600 24124 -416
rect -956 37842 24124 38026
rect -956 -600 -772 38026
rect 23940 -600 24124 38026
rect 24540 -1200 24724 38626
rect -1556 -1200 24724 -1016
rect -1556 38442 24724 38626
rect -1556 -1200 -1372 38626
rect 24540 -1200 24724 38626
rect -1556 39042 24724 39226
rect -1556 39042 24724 39226
rect 24844 -1380 24904 39226
rect -1556 -1380 24904 -1320
rect 24844 -1380 24904 39226
rect -1736 -1560 24904 -1500
rect -1736 -1560 -1676 39226
rect 18514 34116 18694 34176
rect 1354 32756 1534 32816
rect 2734 26996 2914 27056
rect 10774 2450 10954 2510
rect 10774 1170 10954 1230
use SARBSSW_CV XB1
transform -1 0 11584 0 1 0
box 11584 0 23524 4800
use SARBSSW_CV XB2
transform 1 0 11584 0 1 0
box 11584 0 23524 4800
use CDAC8_CV XDAC1
transform -1 0 11404 0 1 4990
box 11404 4990 22692 16954
use CDAC8_CV XDAC2
transform 1 0 11744 0 1 4990
box 11744 4990 23032 16954
use SARDIGEX4_CV XA0
transform 1 0 1084 0 1 23346
box 1084 23346 3184 36466
use SARDIGEX4_CV XA1
transform -1 0 5284 0 1 23346
box 5284 23346 7384 36466
use SARDIGEX4_CV XA2
transform 1 0 5284 0 1 23346
box 5284 23346 7384 36466
use SARDIGEX4_CV XA3
transform -1 0 9484 0 1 23346
box 9484 23346 11584 36466
use SARDIGEX4_CV XA4
transform 1 0 9484 0 1 23346
box 9484 23346 11584 36466
use SARDIGEX4_CV XA5
transform -1 0 13684 0 1 23346
box 13684 23346 15784 36466
use SARDIGEX4_CV XA6
transform 1 0 13684 0 1 23346
box 13684 23346 15784 36466
use SARDIGEX4_CV XA7
transform -1 0 17884 0 1 23346
box 17884 23346 19984 36466
use SARDIGEX4_CV XA8
transform 1 0 17884 0 1 23346
box 17884 23346 19984 36466
use SARCMPX1_CV XA20
transform -1 0 22084 0 1 23346
box 22084 23346 24184 37426
use cut_M3M4_1x2 
transform 1 0 14500 0 1 16954
box 14500 16954 14568 17138
use cut_M3M4_2x1 
transform 1 0 14500 0 1 17456
box 14500 17456 14684 17524
use cut_M3M4_1x2 
transform 1 0 8580 0 1 16954
box 8580 16954 8648 17138
use cut_M3M4_2x1 
transform 1 0 8580 0 1 17836
box 8580 17836 8764 17904
use cut_M2M4_2x1 
transform 1 0 21634 0 1 25396
box 21634 25396 21818 25464
use cut_M4M5_2x1 
transform 1 0 21634 0 1 17836
box 21634 17836 21818 17904
use cut_M4M5_1x2 
transform 1 0 21634 0 1 18176
box 21634 18176 21702 18360
use cut_M3M4_2x1 
transform 1 0 21762 0 1 32436
box 21762 32436 21946 32504
use cut_M2M3_2x1 
transform 1 0 21634 0 1 32436
box 21634 32436 21818 32504
use cut_M4M5_2x1 
transform 1 0 21878 0 1 17456
box 21878 17456 22062 17524
use cut_M4M5_1x2 
transform 1 0 21878 0 1 18176
box 21878 18176 21946 18360
use cut_M3M4_1x2 
transform 1 0 4834 0 1 18158
box 4834 18158 4902 18342
use cut_M2M3_1x2 
transform 1 0 13552 0 1 18158
box 13552 18158 13620 18342
use cut_M3M4_1x2 
transform 1 0 5550 0 1 18348
box 5550 18348 5618 18532
use cut_M2M3_1x2 
transform 1 0 13176 0 1 18348
box 13176 18348 13244 18532
use cut_M3M4_1x2 
transform 1 0 9034 0 1 18538
box 9034 18538 9102 18722
use cut_M2M3_1x2 
transform 1 0 12800 0 1 18538
box 12800 18538 12868 18722
use cut_M3M4_1x2 
transform 1 0 1350 0 1 18728
box 1350 18728 1418 18912
use cut_M2M3_1x2 
transform 1 0 13928 0 1 18728
box 13928 18728 13996 18912
use cut_M3M4_1x2 
transform 1 0 12738 0 1 18918
box 12738 18918 12806 19102
use cut_M2M3_1x2 
transform 1 0 10844 0 1 18918
box 10844 18918 10912 19102
use cut_M3M4_1x2 
transform 1 0 16938 0 1 19108
box 16938 19108 17006 19292
use cut_M2M3_1x2 
transform 1 0 11220 0 1 19108
box 11220 19108 11288 19292
use cut_M3M4_1x2 
transform 1 0 10362 0 1 19298
box 10362 19298 10430 19482
use cut_M2M3_1x2 
transform 1 0 10656 0 1 19298
box 10656 19298 10724 19482
use cut_M3M4_1x2 
transform 1 0 14562 0 1 19488
box 14562 19488 14630 19672
use cut_M2M3_1x2 
transform 1 0 11032 0 1 19488
box 11032 19488 11100 19672
use cut_M3M4_1x2 
transform 1 0 1962 0 1 19678
box 1962 19678 2030 19862
use cut_M2M3_1x2 
transform 1 0 9152 0 1 19678
box 9152 19678 9220 19862
use cut_M3M4_1x2 
transform 1 0 6162 0 1 19868
box 6162 19868 6230 20052
use cut_M2M3_1x2 
transform 1 0 9904 0 1 19868
box 9904 19868 9972 20052
use cut_M3M4_1x2 
transform 1 0 4338 0 1 20058
box 4338 20058 4406 20242
use cut_M2M3_1x2 
transform 1 0 9528 0 1 20058
box 9528 20058 9596 20242
use cut_M3M4_1x2 
transform 1 0 8538 0 1 20248
box 8538 20248 8606 20432
use cut_M2M3_1x2 
transform 1 0 10280 0 1 20248
box 10280 20248 10348 20432
use cut_M3M4_1x2 
transform 1 0 2098 0 1 20438
box 2098 20438 2166 20622
use cut_M2M3_1x2 
transform 1 0 9340 0 1 20438
box 9340 20438 9408 20622
use cut_M3M4_1x2 
transform 1 0 8402 0 1 20628
box 8402 20628 8470 20812
use cut_M2M3_1x2 
transform 1 0 10468 0 1 20628
box 10468 20628 10536 20812
use cut_M3M4_1x2 
transform 1 0 6298 0 1 20818
box 6298 20818 6366 21002
use cut_M2M3_1x2 
transform 1 0 10092 0 1 20818
box 10092 20818 10160 21002
use cut_M3M4_1x2 
transform 1 0 4202 0 1 21008
box 4202 21008 4270 21192
use cut_M2M3_1x2 
transform 1 0 9716 0 1 21008
box 9716 21008 9784 21192
use cut_M3M4_1x2 
transform 1 0 10634 0 1 21198
box 10634 21198 10702 21382
use cut_M2M3_1x2 
transform 1 0 12424 0 1 21198
box 12424 21198 12492 21382
use cut_M3M4_1x2 
transform 1 0 12466 0 1 21388
box 12466 21388 12534 21572
use cut_M2M3_1x2 
transform 1 0 12236 0 1 21388
box 12236 21388 12304 21572
use cut_M3M4_1x2 
transform 1 0 14834 0 1 21578
box 14834 21578 14902 21762
use cut_M2M3_1x2 
transform 1 0 12048 0 1 21578
box 12048 21578 12116 21762
use cut_M3M4_1x2 
transform 1 0 8266 0 1 21768
box 8266 21768 8334 21952
use cut_M2M3_1x2 
transform 1 0 12612 0 1 21768
box 12612 21768 12680 21952
use cut_M3M4_1x2 
transform 1 0 4066 0 1 21958
box 4066 21958 4134 22142
use cut_M2M3_1x2 
transform 1 0 13364 0 1 21958
box 13364 21958 13432 22142
use cut_M3M4_1x2 
transform 1 0 2234 0 1 22148
box 2234 22148 2302 22332
use cut_M2M3_1x2 
transform 1 0 13740 0 1 22148
box 13740 22148 13808 22332
use cut_M3M4_1x2 
transform 1 0 16666 0 1 22338
box 16666 22338 16734 22522
use cut_M2M3_1x2 
transform 1 0 11860 0 1 22338
box 11860 22338 11928 22522
use cut_M3M4_1x2 
transform 1 0 6434 0 1 22528
box 6434 22528 6502 22712
use cut_M2M3_1x2 
transform 1 0 12988 0 1 22528
box 12988 22528 13056 22712
use cut_M1M4_2x2 
transform 1 0 1714 0 1 37842
box 1714 37842 1898 38026
use cut_M1M4_2x2 
transform 1 0 4470 0 1 37842
box 4470 37842 4654 38026
use cut_M1M4_2x2 
transform 1 0 5914 0 1 37842
box 5914 37842 6098 38026
use cut_M1M4_2x2 
transform 1 0 8670 0 1 37842
box 8670 37842 8854 38026
use cut_M1M4_2x2 
transform 1 0 10114 0 1 37842
box 10114 37842 10298 38026
use cut_M1M4_2x2 
transform 1 0 12870 0 1 37842
box 12870 37842 13054 38026
use cut_M1M4_2x2 
transform 1 0 14314 0 1 37842
box 14314 37842 14498 38026
use cut_M1M4_2x2 
transform 1 0 17070 0 1 37842
box 17070 37842 17254 38026
use cut_M1M4_2x2 
transform 1 0 18514 0 1 37842
box 18514 37842 18698 38026
use cut_M1M4_2x2 
transform 1 0 21270 0 1 37842
box 21270 37842 21454 38026
use cut_M1M4_2x2 
transform 1 0 9570 0 1 -600
box 9570 -600 9754 -416
use cut_M1M4_2x2 
transform 1 0 13414 0 1 -600
box 13414 -600 13598 -416
use cut_M1M4_2x2 
transform 1 0 2374 0 1 38442
box 2374 38442 2558 38626
use cut_M1M4_2x2 
transform 1 0 3810 0 1 38442
box 3810 38442 3994 38626
use cut_M1M4_2x2 
transform 1 0 6574 0 1 38442
box 6574 38442 6758 38626
use cut_M1M4_2x2 
transform 1 0 8010 0 1 38442
box 8010 38442 8194 38626
use cut_M1M4_2x2 
transform 1 0 10774 0 1 38442
box 10774 38442 10958 38626
use cut_M1M4_2x2 
transform 1 0 12210 0 1 38442
box 12210 38442 12394 38626
use cut_M1M4_2x2 
transform 1 0 14974 0 1 38442
box 14974 38442 15158 38626
use cut_M1M4_2x2 
transform 1 0 16410 0 1 38442
box 16410 38442 16594 38626
use cut_M1M4_2x2 
transform 1 0 19174 0 1 38442
box 19174 38442 19358 38626
use cut_M1M4_2x2 
transform 1 0 20610 0 1 38442
box 20610 38442 20794 38626
use cut_M1M4_2x2 
transform 1 0 8910 0 1 -1200
box 8910 -1200 9094 -1016
use cut_M1M4_2x2 
transform 1 0 14074 0 1 -1200
box 14074 -1200 14258 -1016
use cut_M1M4_2x2 
transform 1 0 2854 0 1 39042
box 2854 39042 3038 39226
use cut_M1M4_2x2 
transform 1 0 3330 0 1 39042
box 3330 39042 3514 39226
use cut_M1M4_2x2 
transform 1 0 7054 0 1 39042
box 7054 39042 7238 39226
use cut_M1M4_2x2 
transform 1 0 7530 0 1 39042
box 7530 39042 7714 39226
use cut_M1M4_2x2 
transform 1 0 11254 0 1 39042
box 11254 39042 11438 39226
use cut_M1M4_2x2 
transform 1 0 11730 0 1 39042
box 11730 39042 11914 39226
use cut_M1M4_2x2 
transform 1 0 15454 0 1 39042
box 15454 39042 15638 39226
use cut_M1M4_2x2 
transform 1 0 15930 0 1 39042
box 15930 39042 16114 39226
use cut_M1M4_2x2 
transform 1 0 19654 0 1 39042
box 19654 39042 19838 39226
use cut_M1M2_2x1 
transform 1 0 9932 0 1 450
box 9932 450 10116 518
use cut_M1M2_2x1 
transform 1 0 9932 0 1 -1380
box 9932 -1380 10116 -1312
use cut_M1M2_2x1 
transform 1 0 13052 0 1 450
box 13052 450 13236 518
use cut_M1M2_2x1 
transform 1 0 13052 0 1 -1380
box 13052 -1380 13236 -1312
use cut_M1M2_2x1 
transform 1 0 1354 0 1 35636
box 1354 35636 1538 35704
use cut_M1M2_1x2 
transform 1 0 -1740 0 1 35574
box -1740 35574 -1672 35758
use cut_M1M4_2x1 
transform 1 0 10126 0 1 -1560
box 10126 -1560 10310 -1492
use cut_M1M4_2x1 
transform 1 0 12858 0 1 -1560
box 12858 -1560 13042 -1492
use cut_M1M3_2x1 
transform 1 0 2374 0 1 36070
box 2374 36070 2558 36138
use cut_M1M3_2x1 
transform 1 0 4834 0 1 35636
box 4834 35636 5018 35704
use cut_M1M3_2x1 
transform 1 0 6574 0 1 36070
box 6574 36070 6758 36138
use cut_M1M3_2x1 
transform 1 0 9034 0 1 35636
box 9034 35636 9218 35704
use cut_M1M3_2x1 
transform 1 0 10774 0 1 36070
box 10774 36070 10958 36138
use cut_M1M3_2x1 
transform 1 0 13234 0 1 35636
box 13234 35636 13418 35704
use cut_M1M3_2x1 
transform 1 0 14974 0 1 36070
box 14974 36070 15158 36138
use cut_M1M3_2x1 
transform 1 0 17434 0 1 35636
box 17434 35636 17618 35704
use cut_M1M3_2x1 
transform 1 0 1354 0 1 32756
box 1354 32756 1538 32824
use cut_M1M3_2x1 
transform 1 0 4834 0 1 32756
box 4834 32756 5018 32824
use cut_M1M3_2x1 
transform 1 0 5554 0 1 32756
box 5554 32756 5738 32824
use cut_M1M3_2x1 
transform 1 0 9034 0 1 32756
box 9034 32756 9218 32824
use cut_M1M3_2x1 
transform 1 0 9754 0 1 32756
box 9754 32756 9938 32824
use cut_M1M3_2x1 
transform 1 0 13234 0 1 32756
box 13234 32756 13418 32824
use cut_M1M3_2x1 
transform 1 0 13954 0 1 32756
box 13954 32756 14138 32824
use cut_M1M3_2x1 
transform 1 0 17434 0 1 32756
box 17434 32756 17618 32824
use cut_M1M3_2x1 
transform 1 0 18154 0 1 32756
box 18154 32756 18338 32824
use cut_M1M2_2x1 
transform 1 0 3814 0 1 36036
box 3814 36036 3998 36104
use cut_M1M2_2x1 
transform 1 0 5554 0 1 35636
box 5554 35636 5738 35704
use cut_M1M2_2x1 
transform 1 0 8014 0 1 36036
box 8014 36036 8198 36104
use cut_M1M2_2x1 
transform 1 0 9754 0 1 35636
box 9754 35636 9938 35704
use cut_M1M2_2x1 
transform 1 0 12214 0 1 36036
box 12214 36036 12398 36104
use cut_M1M2_2x1 
transform 1 0 13954 0 1 35636
box 13954 35636 14138 35704
use cut_M1M2_2x1 
transform 1 0 16414 0 1 36036
box 16414 36036 16598 36104
use cut_M1M2_2x1 
transform 1 0 18154 0 1 35636
box 18154 35636 18338 35704
use cut_M1M3_2x1 
transform 1 0 1354 0 1 26356
box 1354 26356 1538 26424
use cut_M1M3_2x1 
transform 1 0 4834 0 1 26356
box 4834 26356 5018 26424
use cut_M1M3_2x1 
transform 1 0 5554 0 1 26356
box 5554 26356 5738 26424
use cut_M1M3_2x1 
transform 1 0 9034 0 1 26356
box 9034 26356 9218 26424
use cut_M1M3_2x1 
transform 1 0 9754 0 1 26356
box 9754 26356 9938 26424
use cut_M1M3_2x1 
transform 1 0 13234 0 1 26356
box 13234 26356 13418 26424
use cut_M1M3_2x1 
transform 1 0 13954 0 1 26356
box 13954 26356 14138 26424
use cut_M1M3_2x1 
transform 1 0 17434 0 1 26356
box 17434 26356 17618 26424
use cut_M1M3_2x1 
transform 1 0 18154 0 1 26356
box 18154 26356 18338 26424
use cut_M1M3_2x1 
transform 1 0 2734 0 1 26996
box 2734 26996 2918 27064
use cut_M1M3_2x1 
transform 1 0 2734 0 1 26996
box 2734 26996 2918 27064
use cut_M1M3_2x1 
transform 1 0 3454 0 1 26996
box 3454 26996 3638 27064
use cut_M1M3_2x1 
transform 1 0 6934 0 1 26996
box 6934 26996 7118 27064
use cut_M1M3_2x1 
transform 1 0 7654 0 1 26996
box 7654 26996 7838 27064
use cut_M1M3_2x1 
transform 1 0 11134 0 1 26996
box 11134 26996 11318 27064
use cut_M1M3_2x1 
transform 1 0 11854 0 1 26996
box 11854 26996 12038 27064
use cut_M1M3_2x1 
transform 1 0 15334 0 1 26996
box 15334 26996 15518 27064
use cut_M1M3_2x1 
transform 1 0 16054 0 1 26996
box 16054 26996 16238 27064
use cut_M1M3_2x1 
transform 1 0 19534 0 1 26996
box 19534 26996 19718 27064
use cut_M1M3_2x1 
transform 1 0 21270 0 1 28390
box 21270 28390 21454 28458
use cut_M1M3_2x1 
transform 1 0 20610 0 1 29670
box 20610 29670 20794 29738
use cut_M1M3_2x1 
transform 1 0 20254 0 1 36276
box 20254 36276 20438 36344
use cut_M1M3_2x1 
transform 1 0 18154 0 1 33396
box 18154 33396 18338 33464
use cut_M1M3_2x1 
transform 1 0 20250 0 1 36916
box 20250 36916 20434 36984
use cut_M1M3_2x1 
transform 1 0 19170 0 1 36070
box 19170 36070 19354 36138
use cut_M1M2_2x1 
transform 1 0 20250 0 1 36596
box 20250 36596 20434 36664
use cut_M1M2_2x1 
transform 1 0 18510 0 1 34116
box 18510 34116 18694 34184
use cut_M4M5_1x2 
transform 1 0 10642 0 1 1170
box 10642 1170 10710 1354
use cut_M4M5_1x2 
transform 1 0 10642 0 1 4874
box 10642 4874 10710 5058
use cut_M1M4_2x1 
transform 1 0 12214 0 1 1170
box 12214 1170 12398 1238
use cut_M4M5_1x2 
transform 1 0 12458 0 1 1170
box 12458 1170 12526 1354
use cut_M4M5_1x2 
transform 1 0 12458 0 1 4874
box 12458 4874 12526 5058
use cut_M1M3_2x1 
transform 1 0 10774 0 1 2450
box 10774 2450 10958 2518
use cut_M1M3_2x1 
transform 1 0 12214 0 1 1170
box 12214 1170 12398 1238
use cut_M1M4_2x1 
transform 1 0 10774 0 1 1170
box 10774 1170 10958 1238
use cut_M1M4_2x1 
transform 1 0 12214 0 1 2450
box 12214 2450 12398 2518
use cut_M1M3_2x1 
transform 1 0 1354 0 1 26996
box 1354 26996 1538 27064
use cut_M1M2_2x2 
transform 1 0 -956 0 1 5050
box -956 5050 -772 5234
use cut_M1M2_2x2 
transform 1 0 -956 0 1 6538
box -956 6538 -772 6722
use cut_M1M2_2x2 
transform 1 0 -956 0 1 8026
box -956 8026 -772 8210
use cut_M1M2_2x2 
transform 1 0 -956 0 1 9514
box -956 9514 -772 9698
use cut_M1M2_2x2 
transform 1 0 -956 0 1 11002
box -956 11002 -772 11186
use cut_M1M2_2x2 
transform 1 0 -956 0 1 12490
box -956 12490 -772 12674
use cut_M1M2_2x2 
transform 1 0 -956 0 1 13978
box -956 13978 -772 14162
use cut_M1M2_2x2 
transform 1 0 -956 0 1 15466
box -956 15466 -772 15650
use cut_M1M2_2x2 
transform 1 0 23940 0 1 4990
box 23940 4990 24124 5174
use cut_M1M2_2x2 
transform 1 0 23940 0 1 6478
box 23940 6478 24124 6662
use cut_M1M2_2x2 
transform 1 0 23940 0 1 7966
box 23940 7966 24124 8150
use cut_M1M2_2x2 
transform 1 0 23940 0 1 9454
box 23940 9454 24124 9638
use cut_M1M2_2x2 
transform 1 0 23940 0 1 10942
box 23940 10942 24124 11126
use cut_M1M2_2x2 
transform 1 0 23940 0 1 12430
box 23940 12430 24124 12614
use cut_M1M2_2x2 
transform 1 0 23940 0 1 13918
box 23940 13918 24124 14102
use cut_M1M2_2x2 
transform 1 0 23940 0 1 15406
box 23940 15406 24124 15590
<< labels >>
flabel m3 s 1350 18854 1418 28592 0 FreeSans 400 0 0 0 D<8>
port 1 nsew
flabel m3 s 12738 19044 12806 28614 0 FreeSans 400 0 0 0 D<3>
port 2 nsew
flabel m3 s 16938 19234 17006 28614 0 FreeSans 400 0 0 0 D<1>
port 3 nsew
flabel m3 s 10362 19424 10430 28614 0 FreeSans 400 0 0 0 D<4>
port 4 nsew
flabel m3 s 14562 19614 14630 28614 0 FreeSans 400 0 0 0 D<2>
port 5 nsew
flabel m3 s 6162 19994 6230 28614 0 FreeSans 400 0 0 0 D<6>
port 6 nsew
flabel m3 s 4338 20184 4406 28614 0 FreeSans 400 0 0 0 D<7>
port 7 nsew
flabel m3 s 8538 20374 8606 28614 0 FreeSans 400 0 0 0 D<5>
port 8 nsew
flabel locali s 23940 -600 24124 38026 0 FreeSans 400 0 0 0 AVSS
port 9 nsew
flabel locali s 24540 -1200 24724 38626 0 FreeSans 400 0 0 0 AVDD
port 10 nsew
flabel locali s -1556 39042 24724 39226 0 FreeSans 400 0 0 0 VREF
port 11 nsew
flabel locali s 24844 -1380 24904 39226 0 FreeSans 400 0 0 0 CK_SAMPLE_BSSW
port 12 nsew
flabel locali s 18514 34116 18694 34176 0 FreeSans 400 0 0 0 DONE
port 13 nsew
flabel m3 s 10774 46 10958 114 0 FreeSans 400 0 0 0 SAR_IP
port 14 nsew
flabel m3 s 12210 46 12394 114 0 FreeSans 400 0 0 0 SAR_IN
port 15 nsew
flabel locali s 1354 32756 1534 32816 0 FreeSans 400 0 0 0 CK_SAMPLE
port 16 nsew
flabel locali s 2734 26996 2914 27056 0 FreeSans 400 0 0 0 EN
port 17 nsew
flabel locali s 10774 2450 10954 2510 0 FreeSans 400 0 0 0 SARN
port 18 nsew
flabel locali s 10774 1170 10954 1230 0 FreeSans 400 0 0 0 SARP
port 19 nsew
flabel m3 s 18762 28614 18830 28798 0 FreeSans 400 0 0 0 D<0>
port 20 nsew
<< end >>
